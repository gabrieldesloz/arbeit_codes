
library ieee;
use IEEE.STD_LOGIC_1164.all;
use ieee.math_real.all;
use ieee.numeric_std.all;


entity EJECT_DEAD_TIME is
  port (
    CLK_1us_i   : in  std_logic;  -- 10 MHz / 100 ns maximum resolution                        
    RESET_i 	: in  std_logic;
    PULSE_i     : in  std_logic;  
    PULSE_o    	: out std_logic;
    DEAD_Time_o : out std_logic
    );

end EJECT_DEAD_TIME;


architecture Behavioral of EJECT_DEAD_TIME is

  type FSM_1 is (st_IDLE, st_ACTIVE, st_DEAD_T);
  signal state_reg, state_next               : FSM_1;
   

  constant DEFLUX_T                      : natural := 800;  -- us
  constant MAX_COUNT 				     : natural := DEFLUX_T; 		
  constant DATA_COUNT_bits               : natural := integer(ceil(log2(real(MAX_COUNT))));
  
  signal pulse_i_reg, pulse_i_next: 													    		std_logic; 	
  signal pulse_o_reg, pulse_o_next: 													    		std_logic; 	
  signal dead_time_reg, dead_time_next: 													        std_logic; 	
  signal count_reg, count_next:												            			unsigned(DATA_COUNT_bits-1 downto 0);
  

begin

		
  registers : process (CLK_1us_i, RESET_i)  -- 1MHz
  begin
    
	if (RESET_i = '1') then
	
      state_reg                                   <= st_IDLE;
	  pulse_i_reg								  <= '0';		
	  pulse_o_reg                                 <= '0'; 
	  dead_time_reg                               <= '0';
	  
		
	elsif rising(CLK_1us_i) then
	  
      state_reg                                   <= state_next;
      pulse_i_reg								  <= PULSE_i;		
	  pulse_o_reg                                 <= pulse_o_next;  
	  dead_time_reg                               <= dead_time_next;
	  
    end if;
  end process registers;

   PULSE_o 			<= pulse_o_reg;
   DEAD_Time_o 		<= dead_time_reg;
   
  fsm : process(pulse_i_reg, pulse_o_reg, state_reg, dead_time_reg)

  begin

    --DEFAULT
 
	state_next          <= state_reg;
	pulse_o_next 		<= pulse_o_reg;
	dead_time_next      <= dead_time_reg;
	count_next          <= count_reg;

    case state_reg is

      when st_IDLE =>
                                      
		pulse_o_next 			<= '0';
		
		if pulse_i_reg = '1' then 
			state_next 			<= st_ACTIVE;		
        end if;
	   
	  when st_ACTIVE =>
		
		pulse_o_next 			<= '1';
		
		if pulse_i_reg = '0' then 
		    count_next 			<= (others => '0');
			state_next 			<= st_DEAD_T;
			dead_time_next      <= '1'; 
        end if;
		
	  
	   when st_DEAD_T =>
	   
	    pulse_o_next 			<= '0';
		 
	    if count_reg = DEFLUX_T then 
		   count_next 			<= (others => '0');
		   state_next 			<= st_IDLE;
		   dead_time_next       <= '0' ;     
		else
		   count_next <= count_reg + 1;
        end if;
	 

      when others =>
		state_next <= st_IDLE;

    end case;

  end process fsm;



end Behavioral;



