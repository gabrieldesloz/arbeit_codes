-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'rtl' of entity 'test'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture rtl of test is

begin

end architecture rtl ; -- of test

