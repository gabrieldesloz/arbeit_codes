-------------------------------------------------------------------------------
-- Title      : asbaarda
-- Project    : 
-------------------------------------------------------------------------------
-- File       : teste.vhd
-- Author     :   <s10169@SMKM02>
-- Company    : 
-- Created    : 2014-09-03
-- Last update: 2014-09-03
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2014 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-09-03  1.0      s10169	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity teste is

  generic (
    );

  port (
    );

end teste;

-------------------------------------------------------------------------------

architecture str of teste is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- Component declarations
  -----------------------------------------------------------------------------

begin  -- str

  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

end str;

-------------------------------------------------------------------------------
