-- VHT off
-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /   Vendor: Xilinx
-- \   \   \/    Version: 6.0
--  \   \        Filename: $RCSfile: floating_point_v6_0_unobf.vhd,v $
--  /   /        Date Last Modified: $Date: 2011/06/01 12:58:19 $
-- /___/   /\    Date Created: Dec 2005
-- \   \  /  \
--  \___\/\___\
--
--Device  : All
--Library : xilinxcorelib
--Purpose : Floating-point operator behavioral model
--
--------------------------------------------------------------------------------
-- VHT on
--  (c) Copyright 2005-2009, 2011 Xilinx, Inc. All rights reserved.
--
--  This file contains confidential and proprietary information
--  of Xilinx, Inc. and is protected under U.S. and
--  international copyright and other intellectual property
--  laws.
--
--  DISCLAIMER
--  This disclaimer is not a license and does not grant any
--  rights to the materials distributed herewith. Except as
--  otherwise provided in a valid license issued to you by
--  Xilinx, and to the maximum extent permitted by applicable
--  law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
--  WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
--  AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
--  BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
--  INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
--  (2) Xilinx shall not be liable (whether in contract or tort,
--  including negligence, or under any other theory of
--  liability) for any loss or damage of any kind or nature
--  related to, arising under or in connection with these
--  materials, including for any direct, or any indirect,
--  special, incidental, or consequential loss or damage
--  (including loss of data, profits, goodwill, or any type of
--  loss or damage suffered as a result of any action brought
--  by a third party) even if such damage or loss was
--  reasonably foreseeable or Xilinx had been advised of the
--  possibility of the same.
--
--  CRITICAL APPLICATIONS
--  Xilinx products are not designed or intended to be fail-
--  safe, or for use in any application requiring fail-safe
--  performance, such as life-support or safety devices or
--  systems, Class III medical devices, nuclear facilities,
--  applications related to the deployment of airbags, or any
--  other applications that could lead to death, personal
--  injury, or severe property or environmental damage
--  (individually and collectively, "Critical
--  Applications"). Customer assumes the sole risk and
--  liability of any use of Xilinx products in Critical
--  Applications, subject only to applicable laws and
--  regulations governing limitations on product liability.
--
--  THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
--  PART OF THIS FILE AT ALL TIMES.
--------------------------------------------------------------------------------
-- Generics
--  Constants for generic values are defined in floating_point_v6_0_consts.vhd
--
--  C_XDEVICEFAMILY        : FPGA device family e.g. "virtex6"
--
--  Operators: set the following to: 1 to enable operation
--                                   0 to disable operation (default)
--  C_HAS_ADD              : add operation
--  C_HAS_SUBTRACT         : subtract operation
--  C_HAS_MULTIPLY         : multiply operation
--  C_HAS_DIVIDE           : divide operation
--  C_HAS_SQRT             : squareroot operation
--  C_HAS_COMPARE          : compare operation
--  C_HAS_FIX_TO_FLT       : fixed-point to float-point conversion operation
--  C_HAS_FLT_TO_FIX       : floating-point to fixed-point conversion operation
--  C_HAS_FLT_TO_FLT       : floating-point to floating-point conversion operation
--
--  Precision:
--   Set the following generics to the precision required.
--
--   For fixed-point:
--       iiii.fffff   2's complement scaled binary number,
--                    where i=integer bits, f= fractional bits
--       <-------->   Total bit-width
--            <--->   Fraction bit-width
--   E.g. 64-bit integer C_A_WIDTH = 64, C_A_FRACTION_WIDTH = 0
--
--   For floating-point:
--
--       seeeffffff   s=sign-bit, e=biased exponent, f=fractional part
--       <-------->   Total bit-width
--          1.fffff
--          <----->   Fraction bit-width
--   E.g. single precision C_A_WIDTH = 32, C_A_FRACTION_WIDTH = 24
--        double precision C_A_WIDTH = 64, C_A_FRACTION_WIDTH = 53
--
--  C_A_WIDTH              : Total bit-width of A operand
--  C_A_FRACTION_WIDTH     : Bit-width of fractional part of A operand (inc hidden bit)
--  C_B_WIDTH              : Total bit-width of B operand
--  C_B_FRACTION_WIDTH     : Bit-width of fractional part of B operand (inc hidden bit)
--  C_RESULT_WIDTH         : Total bit-width of result
--  C_RESULT_FRACTION_WIDTH: Bit-width of fractional part of result (inc hidden bit)
--
--  C_COMPARE_OPERATION    : 0 = FLT_PT_UNORDERED             A ? B  unordered i.e. either NaN
--                           1 = FLT_PT_LESS_THAN             A < B
--                           2 = FLT_PT_EQUAL                 A = B
--                           3 = FLT_PRT_LESS_THAN_OR_EQUAL   A <= B
--                           4 = FLT_PT_GREATER_THAN          A > B
--                           5 = FLT_PT_NOT_EQUAL             A <> B
--                           6 = FLT_PT_GREATER_THAN_OR_EQUAL A >= B
--                           7 = FLT_PT_CONDITION_CODE        Flags: m_axis_result_tdata(3 downto 0) == (> , <, =, UN)
--                           8 = FLT_PT_PROGRAMMABLE          Type of comparison specified by OPERATION channel
--
--  C_LATENCY              : Core Latency:
--                           N < 1000 (FLT_PT_MAX_LATENCY)   Latency = N
--                           N = 1000 (FLT_PT_MAX_LATENCY)   Core fully pipelined
--
--  C_OPTIMIZATION         : Architecture optimization:
--                           1 = FLT_PT_SPEED_OPTIMIZED      Optimized for speed
--                           2 = FLT_PT_LOW_LATENCY          Optimized for low-latency
--
--  C_MULT_USAGE           : Level of embedded multiplier (DSP48E1 / DSP48A1) usage:
--                           0 = FLT_PT_NO_USAGE             Logic only, no DSP48s
--                           1 = FLT_PT_MEDIUM_USAGE         Some usage of DSP48s
--                           2 = FLT_PT_FULL_USAGE           Greater usage of DSP48s
--                           3 = FLT_PT_MAX_USAGE            Greatest usage of DSP48s
--
--  C_RATE                 : Maximum number of cycles between inputs
--                           1 = input every cycle
--                           For divide or square-root can set to value higher
--                           to get multi-cycle behavior e.g.
--                           C_A_FRACTION_WIDTH + 1 = serial square-root
--                           C_A_FRACTION_WIDTH + 2 = serial divider
--
--  Exception signals, as defined by IEEE Std 754: set to 1 to provide the exception bit, 0 to omit it
--  C_HAS_UNDERFLOW        : Provide bit in m_axis_result_tuser to indicate when underflow has occurred
--  C_HAS_OVERFLOW         : Provide bit in m_axis_result_tuser to indicate when overflow has occurred
--  C_HAS_INVALID_OP       : Provide bit in m_axis_result_tuser to indicate when invalid operation has been performed
--  C_HAS_DIVIDE_BY_ZERO   : Provide bit in m_axis_result_tuser to indicate when divide-by-zero occurred
--
--  AXI related generics:
--  C_HAS_ACLKEN           : 1 = Provide clock enable input on core, 0 = no clock enable input
--  C_HAS_ARESETN          : 1 = Provide synchronous reset input (active low) on core, 0 = no reset input
--  C_THROTTLE_SCHEME      : Type of AXI handshaking and presence of TREADY signals
--                           1 = Full AXI handshake, use core clock enable to handle backpressure
--                           2 = Full AXI handshake, use output FIFO to handle backpressure
--                           3 = No AXI handshake, no TREADY except inputs when C_RATE > 1
--                           4 = Full AXI handshake on inputs, no TREADY on output
--  C_HAS_A_TUSER          : 1 = A channel has TUSER signal, 0 = no TUSER
--  C_HAS_A_TLAST          : 1 = A channel has TLAST signal, 0 = no TLAST
--  C_HAS_B                : 1 = B channel present (must match operation selection), 0 = no B channel
--  C_HAS_B_TUSER          : 1 = B channel has TUSER signal, 0 = no TUSER
--  C_HAS_B_TLAST          : 1 = B channel has TLAST signal, 0 = no TLAST
--  C_HAS_OPERATION        : 1 = OPERATION channel present (must match operation selection), 0 = no OPERATION channel
--  C_HAS_OPERATION_TUSER  : 1 = OPERATION channel has TUSER signal, 0 = no TUSER
--  C_HAS_OPERATION_TLAST  : 1 = OPERATION channel has TLAST signal, 0 = no TLAST
--  C_HAS_RESULT_TUSER     : 1 = RESULT channel has TUSER signal (any input has TUSER, any exception used), 0 = no TUSER
--  C_HAS_RESULT_TLAST     : 1 = RESULT channel has TLAST signal (any input has TLAST), 0 = no TLAST
--  C_TLAST_RESOLUTION     : Method of generating RESULT channel TLAST signal
--                           1  = use A channel TLAST
--                           2  = use B channel TLAST
--                           3  = use OPERATION channel TLAST
--                           16 = logical OR of TLASTs of all input channels
--                           17 = logical AND of TLASTs of all input channels
--  C_A_TDATA_WIDTH        : Bit width of A TDATA signal: must be C_A_WIDTH rounded up to next byte
--  C_A_TUSER_WIDTH        : Bit width of A TUSER signal (if present): range 1-256
--  C_B_TDATA_WIDTH        : Bit width of B TDATA signal (if present): must be C_A_WIDTH rounded up to next byte
--  C_B_TUSER_WIDTH        : Bit width of B TUSER signal (if present): range 1-256
--  C_OPERATION_TDATA_WIDTH: Bit width of OPERATION TDATA signal (if present): must be 8
--  C_OPERATION_TUSER_WIDTH: Bit width of OPERATION TUSER signal (if present): range 1-256
--  C_RESULT_TDATA_WIDTH   : Bit width of RESULT TDATA signal: must be C_RESULT_WIDTH rounded up to next byte
--  C_RESULT_TUSER_WIDTH   : Bit width of RESULT TUSER signal (if present): must be:
--                           C_A_TUSER_WIDTH (if C_HAS_A_TUSER) +
--                           C_B_TUSER_WIDTH (if C_HAS_B_TUSER) +
--                           C_OPERATION_TUSER_WIDTH (if C_HAS_OPERATION_TUSER) +
--                           1 for each exception bit provided
--
-- Ports
--  Global inputs:
--   aclk                  : Clock (all signals are synchronous to rising edge of clock)
--   aclken                : enables clock on all registers
--   aresetn               : synchronous reset, active LOW (only resets control, not datapath)
--  AXI channels:            Each channel has TVALID, TREADY (optional), TDATA, TUSER (optional) and TLAST (optional).
--   a                     : AXI4-Stream slave channel for operand A (fixed or floating point)
--   b                     : AXI4-Stream slave channel for operand B (floating point)
--   operation             : AXI4-Stream slave channel for operation control:
--                           (   7   6    5   4   3    2   1   0  )  s_axis_operation_tdata
--                            <-unused-><-cmp_mode--><--prim_op-->
--                           std_logic_vector constants for values are defined in floating_point_v6_0_consts.vhd.
--                           Primary Operation Code (prim_op)
--                            "000" = FLT_PT_ADD_OP_CODE_SLV            Add
--                            "001" = FLT_PT_SUBTRACT_OP_CODE_SLV       Subtract
--                            "100" = FLT_PT_COMPARE_OP_CODE_SLV        Compare
--                            All other values are reserved.
--                           Compare Operation Code (cmp_op) when prim_op is "100" = FLT_PT_COMPARE_OP_CODE_SLV:
--                            "000" = FLT_PT_UNORDERED_SLV              A ? B  (A or B is NaN)
--                            "001" = FLT_PT_LESS_THAN_SLV              A < B
--                            "010" = FLT_PT_EQUAL_SLV                  A = B
--                            "011" = FLT_PRT_LESS_THAN_OR_EQUAL_SLV    A <= B
--                            "100" = FLT_PT_GREATER_THAN_SLV           A > B
--                            "101" = FLT_PT_NOT_EQUAL_SLV              A <> B
--                            "110" = FLT_PT_GREATER_THAN_OR_EQUAL_SLV  A >= B
--                            All other values are reserved.
--   result                : Result of operation (fixed or floating point, or comparison result or condition code)
--                           Exception bits are in TUSER LSBs: from bit 0 upwards:
--                           UNDERFLOW, OVERFLOW, INVALID OPERATION, DIVIDE BY ZERO (each present only if requested)
--------------------------------------------------------------------------------

LIBRARY IEEE;USE IEEE.STD_LOGIC_1164.ALL;USE IEEE.NUMERIC_STD.ALL;USE IEEE.MATH_REAL.ALL;LIBRARY XILINXCORELIB;USE XILINXCORELIB.
BIP_UTILS_PKG_V2_0.ALL;USE XILINXCORELIB.AXI_UTILS_PKG_V1_1.ALL;USE XILINXCORELIB.AXI_UTILS_V1_1_COMPS.ALL;USE XILINXCORELIB.
FLOATING_POINT_V6_0_CONSTS.ALL;USE XILINXCORELIB.FLOATING_POINT_PKG_V6_0.ALL;ENTITY FLOATING_POINT_V6_0 IS GENERIC(C_XDEVICEFAMILY:
STRING:="no_family";C_HAS_ADD:INTEGER:=1;C_HAS_SUBTRACT:INTEGER:=0;C_HAS_MULTIPLY:INTEGER:=0;C_HAS_DIVIDE:INTEGER:=0;C_HAS_SQRT:
INTEGER:=0;C_HAS_COMPARE:INTEGER:=0;C_HAS_FIX_TO_FLT:INTEGER:=0;C_HAS_FLT_TO_FIX:INTEGER:=0;C_HAS_FLT_TO_FLT:INTEGER:=0;C_HAS_RECIP
:INTEGER:=0;C_HAS_RECIP_SQRT:INTEGER:=0;C_A_WIDTH:INTEGER:=32;C_A_FRACTION_WIDTH:INTEGER:=24;C_B_WIDTH:INTEGER:=32;
C_B_FRACTION_WIDTH:INTEGER:=24;C_RESULT_WIDTH:INTEGER:=32;C_RESULT_FRACTION_WIDTH:INTEGER:=24;C_COMPARE_OPERATION:INTEGER:=1;
C_LATENCY:INTEGER:=1000;C_OPTIMIZATION:INTEGER:=1;C_MULT_USAGE:INTEGER:=2;C_RATE:INTEGER:=1;C_HAS_UNDERFLOW:INTEGER:=0;
C_HAS_OVERFLOW:INTEGER:=0;C_HAS_INVALID_OP:INTEGER:=0;C_HAS_DIVIDE_BY_ZERO:INTEGER:=0;C_HAS_ACLKEN:INTEGER:=0;C_HAS_ARESETN:INTEGER
:=0;C_THROTTLE_SCHEME:INTEGER:=1;C_HAS_A_TUSER:INTEGER:=0;C_HAS_A_TLAST:INTEGER:=0;C_HAS_B:INTEGER:=1;C_HAS_B_TUSER:INTEGER:=0;
C_HAS_B_TLAST:INTEGER:=0;C_HAS_OPERATION:INTEGER:=0;C_HAS_OPERATION_TUSER:INTEGER:=0;C_HAS_OPERATION_TLAST:INTEGER:=0;
C_HAS_RESULT_TUSER:INTEGER:=0;C_HAS_RESULT_TLAST:INTEGER:=0;C_TLAST_RESOLUTION:INTEGER:=1;C_A_TDATA_WIDTH:INTEGER:=32;
C_A_TUSER_WIDTH:INTEGER:=1;C_B_TDATA_WIDTH:INTEGER:=32;C_B_TUSER_WIDTH:INTEGER:=1;C_OPERATION_TDATA_WIDTH:INTEGER:=8;
C_OPERATION_TUSER_WIDTH:INTEGER:=1;C_RESULT_TDATA_WIDTH:INTEGER:=32;C_RESULT_TUSER_WIDTH:INTEGER:=1);PORT(ACLK:IN STD_LOGIC:='0';
ACLKEN:IN STD_LOGIC:='1';ARESETN:IN STD_LOGIC:='1';S_AXIS_A_TVALID:IN STD_LOGIC:='0';S_AXIS_A_TREADY:OUT STD_LOGIC:='0';
S_AXIS_A_TDATA:IN STD_LOGIC_VECTOR(C_A_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');S_AXIS_A_TUSER:IN STD_LOGIC_VECTOR(C_A_TUSER_WIDTH-1
 DOWNTO 0):=(OTHERS=>'0');S_AXIS_A_TLAST:IN STD_LOGIC:='0';S_AXIS_B_TVALID:IN STD_LOGIC:='0';S_AXIS_B_TREADY:OUT STD_LOGIC:='0';
S_AXIS_B_TDATA:IN STD_LOGIC_VECTOR(C_B_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');S_AXIS_B_TUSER:IN STD_LOGIC_VECTOR(C_B_TUSER_WIDTH-1
 DOWNTO 0):=(OTHERS=>'0');S_AXIS_B_TLAST:IN STD_LOGIC:='0';S_AXIS_OPERATION_TVALID:IN STD_LOGIC:='0';S_AXIS_OPERATION_TREADY:OUT
 STD_LOGIC:='0';S_AXIS_OPERATION_TDATA:IN STD_LOGIC_VECTOR(C_OPERATION_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');S_AXIS_OPERATION_TUSER
:IN STD_LOGIC_VECTOR(C_OPERATION_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');S_AXIS_OPERATION_TLAST:IN STD_LOGIC:='0';
M_AXIS_RESULT_TVALID:OUT STD_LOGIC:='0';M_AXIS_RESULT_TREADY:IN STD_LOGIC:='0';M_AXIS_RESULT_TDATA:OUT STD_LOGIC_VECTOR(
C_RESULT_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');M_AXIS_RESULT_TUSER:OUT STD_LOGIC_VECTOR(C_RESULT_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS
=>'0');M_AXIS_RESULT_TLAST:OUT STD_LOGIC:='0');END;ARCHITECTURE BEHAVIORAL OF FLOATING_POINT_V6_0 IS FUNCTION
 II1IOOO1II0l1lOl00I1O001I00O0IIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII,IOO0111OO0lOOl10l1l000l0OlI0IIIIII:INTEGER;IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII:STD_LOGIC_VECTOR)RETURN BOOLEAN IS VARIABLE IOOOlI0llOIl11IO01100OI1llOIIOIIII:STD_LOGIC_VECTOR(IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII'length-1 DOWNTO 0
);VARIABLE IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII:STD_LOGIC_VECTOR(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-1 DOWNTO 0);BEGIN IOOOlI0llOIl11IO01100OI1llOIIOIIII:=IIlO1lIIlOlOOO0l10OI1ll0I0O10IIIII;IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII:=IOOOlI0llOIl11IO01100OI1llOIIOIIII(IOOOlI0llOIl11IO01100OI1llOIIOIIII'left DOWNTO IOOOlI0llOIl11IO01100OI1llOIIOIIII'left-IO1lll0I0l0l1ll1O01Ol0III011IOIIII+1);RETURN(IO1IOOl1111OI1OOII1IOl0lIIIIOIIIII(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-2 DOWNTO IOO0111OO0lOOl10l1l000l0OlI0IIIIII
-1)=FLT_PT_ZERO(IO1lll0I0l0l1ll1O01Ol0III011IOIIII-IOO0111OO0lOOl10l1l000l0OlI0IIIIII-1 DOWNTO 0));END;FUNCTION II1001IO0010Oll1I01lOI0I0IlIOIIIII(IO110I1O0010OIOlIO00l1IIOl0llIIIII:SIGNED;IIIOOIO01011011IOIIlllIIOO0l1IIIII:NATURAL)RETURN SIGNED IS VARIABLE II1IOOO00I0OI0O01I000O100llOOIIIII:SIGNED(IO110I1O0010OIOlIO00l1IIOl0llIIIII'range):=IO110I1O0010OIOlIO00l1IIOl0llIIIII;
BEGIN FOR II00OI0110lI1II101lO1OO00I10OIIIII IN 1 TO IIIOOIO01011011IOIIlllIIOO0l1IIIII LOOP II1IOOO00I0OI0O01I000O100llOOIIIII:=II1IOOO00I0OI0O01I000O100llOOIIIII(II1IOOO00I0OI0O01I000O100llOOIIIII'left)&II1IOOO00I0OI0O01I000O100llOOIIIII(II1IOOO00I0OI0O01I000O100llOOIIIII'left DOWNTO II1IOOO00I0OI0O01I000O100llOOIIIII'right+1);END LOOP;RETURN II1IOOO00I0OI0O01I000O100llOOIIIII;END;FUNCTION
 II00OIlIlO101I0IIOO0O1I0ll0OIIIIII(IOOI1l1OO01O111lO010OlO1O0l0IIIIII:UNSIGNED;IO11OllII1lO110Ol0I0O00I01l00IIIII:NATURAL)RETURN UNSIGNED IS VARIABLE III01lO1l00IOOO0O0I0O0I111O0IIIIII:UNSIGNED(IOOI1l1OO01O111lO010OlO1O0l0IIIIII'range):=IOOI1l1OO01O111lO010OlO1O0l0IIIIII;BEGIN FOR IO1I1l01l1OI111Ol0IO10110I11IOIIII IN 1 TO IO11OllII1lO110Ol0I0O00I01l00IIIII LOOP III01lO1l00IOOO0O0I0O0I111O0IIIIII:='0'&
III01lO1l00IOOO0O0I0O0I111O0IIIIII(III01lO1l00IOOO0O0I0O0I111O0IIIIII'left DOWNTO III01lO1l00IOOO0O0I0O0I111O0IIIIII'right+1);END LOOP;RETURN III01lO1l00IOOO0O0I0O0I111O0IIIIII;END;PROCEDURE IOOll1I1OOlO0lOO0IIII1lO11IIlIIIII(IIIOI11O0OO00OllOllO00lOI000IOIIII:IN INTEGER;IIOIOOO11l0lO001OI10I0IIIIlIIIIIII:IN INTEGER;II0IO0I0Olll01OOO0lIOO01lOlIOOIIII:IN
 STD_LOGIC_VECTOR;IOO10IlOOIIIlOIO1IOI1l1lOIIlOIIIII:OUT STD_LOGIC_VECTOR;II0l0OlOIIIO1I0IOlIIllOIOO10lIIIII:OUT STD_LOGIC;IO0lIOlI0II1000IOlOIlOI1lIlOOIIIII:OUT STD_LOGIC;IO0O10O101OOIOOl10lIIO101lIIIIIIII:OUT STD_LOGIC)IS CONSTANT IIOl10001I1Ol001OIO01IO1II10OIIIII:
INTEGER:=IIOIOOO11l0lO001OI10I0IIIIlIIIIIII;CONSTANT IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII:INTEGER:=IIIOI11O0OO00OllOllO00lOI000IOIIII-IIOIOOO11l0lO001OI10I0IIIIlIIIIIII;CONSTANT IIIIl1100lOI0I1OO1I00OlI0l10IIIIII:INTEGER:=2**(IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-1)-1;CONSTANT IOlI00I100IOOOl011O11IOI1l010IIIII:INTEGER:=2-2**(IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-1);CONSTANT
 IIIO1O1110Oll10OI110OIIO111OOIIIII:INTEGER:=2**(IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-1)-1;VARIABLE IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:STD_LOGIC_VECTOR(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 0);VARIABLE IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:STD_LOGIC_VECTOR(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-1 DOWNTO 0);
VARIABLE II11I0011I0IIIl0100l1O01O01O0IIIII:STD_LOGIC:='0';VARIABLE II011lO0O1l10O0I0OIOO000I0O1IOIIII:SIGNED(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 0);VARIABLE IO1IIIl1OO00II0ll110l0l0IIO0lIIIII:INTEGER;VARIABLE IIlOllOOI0ll11O1101IIl0l11ll1IIIII:STD_LOGIC;VARIABLE
 II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:STD_LOGIC_VECTOR(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 0);VARIABLE III1OO10l11110IO1IO0lOII0OO11IIIII:STD_LOGIC;VARIABLE IO1O1llOO0IlllI1O1OlOI010l1IIIIIII:INTEGER;VARIABLE IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:SIGNED(IIOl10001I1Ol001OIO01IO1II10OIIIII+3 DOWNTO 0);BEGIN
 II11I0011I0IIIl0100l1O01O01O0IIIII:='0';IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:=(OTHERS=>'0');IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:=(OTHERS=>'0');IIlOllOOI0ll11O1101IIl0l11ll1IIIII:=II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-1);IF FLT_PT_IS_NAN(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII,II0IO0I0Olll01OOO0lIOO01lOlIOOIIII)THEN IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=FLT_PT_GET_QUIET_NAN(
IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII);ELSIF II1IOOO1II0l1lOl00I1O001I00O0IIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII,II0IO0I0Olll01OOO0lIOO01lOlIOOIIII)THEN IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=FLT_PT_GET_ZERO(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII,IIlOllOOI0ll11O1101IIl0l11ll1IIIII);ELSIF IIlOllOOI0ll11O1101IIl0l11ll1IIIII='1'THEN II11I0011I0IIIl0100l1O01O01O0IIIII:='1';
IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=FLT_PT_GET_QUIET_NAN(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII);ELSIF FLT_PT_IS_INF(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII,II0IO0I0Olll01OOO0lIOO01lOlIOOIIII)THEN IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=FLT_PT_GET_INF(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII,IIOl10001I1Ol001OIO01IO1II10OIIIII,IIlOllOOI0ll11O1101IIl0l11ll1IIIII);ELSE II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII):=
'1';II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII-1 DOWNTO 1):=SIGNED(II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII-2 DOWNTO 0));II011lO0O1l10O0I0OIOO000I0O1IOIIII(0):='0';IO1IIIl1OO00II0ll110l0l0IIO0lIIIII:=TO_INTEGER(UNSIGNED(II0IO0I0Olll01OOO0lIOO01lOlIOOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII+IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII-2 DOWNTO IIOl10001I1Ol001OIO01IO1II10OIIIII-1)));IF IIlOllOOI0ll11O1101IIl0l11ll1IIIII='1'
THEN III1OO10l11110IO1IO0lOII0OO11IIIII:='1';ELSE III1OO10l11110IO1IO0lOII0OO11IIIII:='0';END IF;IO1O1llOO0IlllI1O1OlOI010l1IIIIIII:=(IO1IIIl1OO00II0ll110l0l0IIO0lIIIII+IIIIl1100lOI0I1OO1I00OlI0l10IIIIII)/2;IF(IO1IIIl1OO00II0ll110l0l0IIO0lIIIII MOD 2=1)THEN II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 0):='0'&II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII
 DOWNTO 1);END IF;FOR II1IO01lI1IO1OII11O1II01I0llIOIIII IN(IIOl10001I1Ol001OIO01IO1II10OIIIII)DOWNTO 0 LOOP IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:=IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII+1 DOWNTO 0)&SIGNED(II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO IIOl10001I1Ol001OIO01IO1II10OIIIII-1));IF IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII>=0 THEN IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:=IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII-SIGNED(RESIZE(
UNSIGNED(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII&"01"),IIOl10001I1Ol001OIO01IO1II10OIIIII+3));ELSE IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII:=IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII+SIGNED(RESIZE(UNSIGNED(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII&"11"),IIOl10001I1Ol001OIO01IO1II10OIIIII+3));END IF;IF IO1O0llO0I1lI11I1O10I0l1O0l0IIIIII>=0 THEN IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:=IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII-1 DOWNTO 0)&'1';ELSE IIl0OIlO00I0lI101l1I0lO1II0IlIIIII:=IIl0OIlO00I0lI101l1I0lO1II0IlIIIII
(IIOl10001I1Ol001OIO01IO1II10OIIIII-1 DOWNTO 0)&'0';END IF;II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 0):=II011lO0O1l10O0I0OIOO000I0O1IOIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII-2 DOWNTO 0)&"00";END LOOP;IF(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(0)='1')THEN II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=STD_LOGIC_VECTOR(
RESIZE(UNSIGNED(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 1)),IIOl10001I1Ol001OIO01IO1II10OIIIII+1)+1);ELSE II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IIl0OIlO00I0lI101l1I0lO1II0IlIIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII DOWNTO 1)),IIOl10001I1Ol001OIO01IO1II10OIIIII+1));END IF;IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII:=
III1OO10l11110IO1IO0lOII0OO11IIIII&STD_LOGIC_VECTOR(TO_UNSIGNED(IO1O1llOO0IlllI1O1OlOI010l1IIIIIII,IIIO0lOII1OIlOOIO1IlI1lIIO001IIIII))&II1I0lOOIIOI1l0l10l0O0l0Ol0OIIIIII(IIOl10001I1Ol001OIO01IO1II10OIIIII-2 DOWNTO 0);END IF;IOO10IlOOIIIlOIO1IOI1l1lOIIlOIIIII:=IOIlII1I0O0l1l1O110O0IOlO0O1lIIIII;II0l0OlOIIIO1I0IOlIIllOIOO10lIIIII:=II11I0011I0IIIl0100l1O01O01O0IIIII;IO0lIOlI0II1000IOlOIlOI1lIlOOIIIII:='0';
IO0O10O101OOIOOl10lIIO101lIIIIIIII:='0';END;PROCEDURE II1lIII001001Il0l0OOl0I00I01IIIIII(II0O0l0l00OIOl0Ol101Il1Ol0I1lIIIII:IN INTEGER;IOII100I0I1l010IOI1lO1O1I1101IIIII:IN INTEGER;IOO10OI11Il110I11IIIIIOIO10OlIIIII:IN STD_LOGIC_VECTOR;IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII:IN STD_LOGIC_VECTOR;IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:OUT
 STD_LOGIC_VECTOR;IOO1l1010O10O10I0llO11O100O1IOIIII:OUT STD_LOGIC;IOIlOIOl1lO1l001Ol10IO01OIlI1IIIII:OUT STD_LOGIC;II0IOOI1Il101lO1O010O0O0IO10IOIIII:OUT STD_LOGIC;IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII:OUT STD_LOGIC)IS CONSTANT
 IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII:INTEGER:=IOII100I0I1l010IOI1lO1O1I1101IIIII;CONSTANT II111OIOII1IIOOOlO1I011OI0I0lIIIII:INTEGER:=II0O0l0l00OIOl0Ol101Il1Ol0I1lIIIII-IOII100I0I1l010IOI1lO1O1I1101IIIII;CONSTANT III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII:INTEGER:=2**(II111OIOII1IIOOOlO1I011OI0I0lIIIII-1)-1;CONSTANT IIIIlI10IO0IlIll11O0O1OII0OIIOIIII:INTEGER:=2-2**(II111OIOII1IIOOOlO1I011OI0I0lIIIII-1);CONSTANT
 IIIO10O1ll1l0O0IOl0l1lllO0lI1IIIII:INTEGER:=2**(II111OIOII1IIOOOlO1I011OI0I0lIIIII-1)-1;VARIABLE IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII:STD_LOGIC_VECTOR(II111OIOII1IIOOOlO1I011OI0I0lIIIII+1 DOWNTO 0);VARIABLE IIl1O1I0001l1001OllOOII0I10l1IIIII:STD_LOGIC_VECTOR(II111OIOII1IIOOOlO1I011OI0I0lIIIII+1 DOWNTO 0);VARIABLE
 IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:SIGNED(II111OIOII1IIOOOlO1I011OI0I0lIIIII+1 DOWNTO 0);VARIABLE IOOI10l0O1lIlIll00Ol1lll10IIIIIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0);VARIABLE IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0);VARIABLE
 IOl0I10010lIIIl000I1O1IO1IlOIIIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0);VARIABLE IOl1I1O0IIO001llOlll1I1lOI1l0IIIII:STD_LOGIC;VARIABLE IOl1Ol11IlIl0110l0OOll000lI11IIIII:STD_LOGIC;VARIABLE II001Il0III1O1OI001IOI100000OIIIII:STD_LOGIC;VARIABLE IOOl0llO0OI110111OIOlOIO0lOOIOIIII:
BOOLEAN;VARIABLE II1IOO1l1I11I1ll1OI1I00lII000IIIII:BOOLEAN;VARIABLE II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII:BOOLEAN;VARIABLE IOOl0IOOO1011llOIOl01lIOI0O11IIIII:BOOLEAN;VARIABLE IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII:BOOLEAN;VARIABLE II1I0O0100lIIII11lI00l0OOII0lIIIII:BOOLEAN;CONSTANT IIOIOI0lO1lO100O11Il0OII11OlOIIIII
:INTEGER:=2;VARIABLE IO0IlO1lI10Il011101l101IIl0IOIIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII-1 DOWNTO 0);VARIABLE IOI1O00I10101l0I1001llOOI0I0IOIIII:STD_LOGIC;VARIABLE IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:STD_LOGIC;
VARIABLE IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:STD_LOGIC;VARIABLE IO0l0IOllOl1100O10O1O1l0lIO1OIIIII:STD_LOGIC;VARIABLE IIlOO000I01110Ill0l1OI1l10IOIOIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1+IIOIOI0lO1lO100O11Il0OII11OlOIIIII+1 DOWNTO 0);VARIABLE II1011O1IO1l0llOI11lIIOIlOlIlIIIII:
UNSIGNED(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0);VARIABLE IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:SIGNED(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO 0);VARIABLE IOI01l1I0000lIO0IIO01IlIO1001IIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO 0);VARIABLE IOI0IIll0I0l1IO0I01lO110IIIIIOIIII:STD_LOGIC;
VARIABLE IO00l1I0I1IOlII011Il0l0lOI0OIIIIII:STD_LOGIC;VARIABLE IO01l1ll0IlOll0I00lll11l0OllIIIIII:STD_LOGIC;VARIABLE IOI11IOIlOI1II1Il11OlI01Illl0IIIII:STD_LOGIC_VECTOR(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO 0);VARIABLE IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII:UNSIGNED(0 DOWNTO 0);
VARIABLE IOlIOOI0O1OIlOl01O0OIII10O11lIIIII:STD_LOGIC;BEGIN IOI1O00I10101l0I1001llOOI0I0IOIIII:='0';IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:='0';IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:='0';IO0l0IOllOl1100O10O1O1l0lIO1OIIIII:='0';IOl1I1O0IIO001llOlll1I1lOI1l0IIIII:=IOO10OI11Il110I11IIIIIOIO10OlIIIII(II111OIOII1IIOOOlO1I011OI0I0lIIIII+IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1);IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII
:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IOO10OI11Il110I11IIIIIOIO10OlIIIII(II111OIOII1IIOOOlO1I011OI0I0lIIIII+IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-2 DOWNTO IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1)),II111OIOII1IIOOOlO1I011OI0I0lIIIII+2));IOOI10l0O1lIlIll00Ol1lll10IIIIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0):='1'&IOO10OI11Il110I11IIIIIOIO10OlIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-2 DOWNTO 0);IOl1Ol11IlIl0110l0OOll000lI11IIIII:=IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII(II111OIOII1IIOOOlO1I011OI0I0lIIIII+IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1);IIl1O1I0001l1001OllOOII0I10l1IIIII
:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII(II111OIOII1IIOOOlO1I011OI0I0lIIIII+IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-2 DOWNTO IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1)),II111OIOII1IIOOOlO1I011OI0I0lIIIII+2));IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0):='1'&IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-2 DOWNTO 0);II001Il0III1O1OI001IOI100000OIIIII:=(IOl1I1O0IIO001llOlll1I1lOI1l0IIIII XOR IOl1Ol11IlIl0110l0OOll000lI11IIIII
);IOOl0llO0OI110111OIOlOIO0lOOIOIIII:=FLT_PT_IS_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO10OI11Il110I11IIIIIOIO10OlIIIII);II1IOO1l1I11I1ll1OI1I00lII000IIIII:=FLT_PT_IS_NAN(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO10OI11Il110I11IIIIIOIO10OlIIIII);II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO10OI11Il110I11IIIIIOIO10OlIIIII);IOOl0IOOO1011llOIOl01lIOI0O11IIIII:=FLT_PT_IS_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII
+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII);IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII:=FLT_PT_IS_NAN(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII);II1I0O0100lIIII11lI00l0OOII0lIIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,IOO1I1lI11Ol1l1OOlllIIII1l1IOIIIII);IF(II1IOO1l1I11I1ll1OI1I00lII000IIIII OR IIOlOO00Ol0011IIIIIO1I1lllIO0IIIII)THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_QUIET_NAN(
IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII);ELSIF IOOl0llO0OI110111OIOlOIO0lOOIOIIII THEN IF IOOl0IOOO1011llOIOl01lIOI0O11IIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_QUIET_NAN(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII:='1';ELSIF II1I0O0100lIIII11lI00l0OOII0lIIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII
,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);ELSE IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);END IF;ELSIF II0II1IO1I0IOIl0ll1I0O00lIIOOIIIII THEN IF IOOl0IOOO1011llOIOl01lIOI0O11IIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_ZERO(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);ELSIF
 II1I0O0100lIIII11lI00l0OOII0lIIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_QUIET_NAN(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII);IOI1O00I10101l0I1001llOOI0I0IOIIII:='1';ELSE IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_ZERO(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);END IF;ELSE IF IOOl0IOOO1011llOIOl01lIOI0O11IIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII
:=FLT_PT_GET_ZERO(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);ELSIF II1I0O0100lIIII11lI00l0OOII0lIIIII THEN IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=FLT_PT_GET_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);IO0l0IOllOl1100O10O1O1l0lIO1OIIIII:='1';ELSE IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:=SIGNED(IIIlOO0OOl101Ol0Oll10O1lOIIO0IIIII)-
SIGNED(IIl1O1I0001l1001OllOOII0I10l1IIIII);IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0):=SIGNED(IOOI10l0O1lIlIll00Ol1lll10IIIIIIII);IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII):=(OTHERS=>'0');IOI01l1I0000lIO0IIO01IlIO1001IIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1 DOWNTO 0):=IO0OOOI1IIIlIOIIOO0Il00I1lOOlIIIII;IOI01l1I0000lIO0IIO01IlIO1001IIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII):=(
OTHERS=>'0');FOR IO1OIOI0I1l11O0IllIOllII1llIIOIIII IN IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+IIOIOI0lO1lO100O11Il0OII11OlOIIIII DOWNTO 1 LOOP IF IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1)='0'THEN IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:=IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII-SIGNED(IOI01l1I0000lIO0IIO01IlIO1001IIIII);IIlOO000I01110Ill0l1OI1l10IOIOIIII(IO1OIOI0I1l11O0IllIOllII1llIIOIIII):='1';ELSE IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:=IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII+SIGNED(IOI01l1I0000lIO0IIO01IlIO1001IIIII);IIlOO000I01110Ill0l1OI1l10IOIOIIII(IO1OIOI0I1l11O0IllIOllII1llIIOIIII):='0';
END IF;IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1 DOWNTO 1):=IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII DOWNTO 0);IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(0):='0';END LOOP;IF IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+1)='0'THEN IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:=IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII-SIGNED(IOI01l1I0000lIO0IIO01IlIO1001IIIII);IIlOO000I01110Ill0l1OI1l10IOIOIIII(0):='1';ELSE IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII:=IOO0I1l1IOO0II0O00I0IllOOI1OOIIIII
+SIGNED(IOI01l1I0000lIO0IIO01IlIO1001IIIII);IIlOO000I01110Ill0l1OI1l10IOIOIIII(0):='0';END IF;IIlOO000I01110Ill0l1OI1l10IOIOIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+IIOIOI0lO1lO100O11Il0OII11OlOIIIII DOWNTO 0):=IIlOO000I01110Ill0l1OI1l10IOIOIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-1+IIOIOI0lO1lO100O11Il0OII11OlOIIIII DOWNTO 0)&'1';IOI0IIll0I0l1IO0I01lO110IIIIIOIIII:=IIlOO000I01110Ill0l1OI1l10IOIOIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+IIOIOI0lO1lO100O11Il0OII11OlOIIIII);IF(IOI0IIll0I0l1IO0I01lO110IIIIIOIIII='1')THEN IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII(0):=IIlOO000I01110Ill0l1OI1l10IOIOIIII(IIOIOI0lO1lO100O11Il0OII11OlOIIIII);II1011O1IO1l0llOI11lIIOIlOlIlIIIII
:=UNSIGNED(IIlOO000I01110Ill0l1OI1l10IOIOIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+IIOIOI0lO1lO100O11Il0OII11OlOIIIII DOWNTO IIOIOI0lO1lO100O11Il0OII11OlOIIIII+1))+IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII;ELSE IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII-1;IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII(0):=IIlOO000I01110Ill0l1OI1l10IOIOIIII(IIOIOI0lO1lO100O11Il0OII11OlOIIIII-1);II1011O1IO1l0llOI11lIIOIlOlIlIIIII:=UNSIGNED(IIlOO000I01110Ill0l1OI1l10IOIOIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+IIOIOI0lO1lO100O11Il0OII11OlOIIIII-1 DOWNTO IIOIOI0lO1lO100O11Il0OII11OlOIIIII))+IIlO0IOl0I0I0lI0OOll1l1l1lO0IIIIII;END IF
;IF TO_INTEGER(IIlIlll0III10I0Il0I0OOOIOIIOOIIIII)>IIIO10O1ll1l0O0IOl0l1lllO0lI1IIIII THEN IO0IlO1lI10Il011101l101IIl0IOIIIII:=FLT_PT_GET_INF(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII:='1';ELSIF TO_INTEGER(IIlIlll0III10I0Il0I0OOOIOIIOOIIIII)<IIIIlI10IO0IlIll11O0O1OII0OIIOIIII THEN
 IO0IlO1lI10Il011101l101IIl0IOIIIII:=FLT_PT_GET_ZERO(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII+II111OIOII1IIOOOlO1I011OI0I0lIIIII,IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII,II001Il0III1O1OI001IOI100000OIIIII);IO1Il1I0OOOOIl0IOO011l1I0111OIIIII:='1';ELSE IIlIlll0III10I0Il0I0OOOIOIIOOIIIII:=IIlIlll0III10I0Il0I0OOOIOIIOOIIIII+III0OI0OlIOOl1Ol1I0l00O0lI1IIIIIII;IO0IlO1lI10Il011101l101IIl0IOIIIII:=II001Il0III1O1OI001IOI100000OIIIII&STD_LOGIC_VECTOR(IIlIlll0III10I0Il0I0OOOIOIIOOIIIII(II111OIOII1IIOOOlO1I011OI0I0lIIIII-1
 DOWNTO 0))&STD_LOGIC_VECTOR(II1011O1IO1l0llOI11lIIOIlOlIlIIIII(IOOIOOI00l1OOOlI1OOO0I00Ol0IlIIIII-2 DOWNTO 0));END IF;IOl0l10lI11IO10lI1OI1IOI01OO0IIIII:=IO0IlO1lI10Il011101l101IIl0IOIIIII;END IF;END IF;IOO1l1010O10O10I0llO11O100O1IOIIII:=IOI1O00I10101l0I1001llOOI0I0IOIIII;IO1lIIIOl1IIIO1O1lllOO0I1lO0OIIIII:=
IO0l0IOllOl1100O10O1O1l0lIO1OIIIII;IOIlOIOl1lO1l001Ol10IO01OIlI1IIIII:=IIOIO000I1OI0OlOI1OIOI1l0I0l1IIIII;II0IOOI1Il101lO1O010O0O0IO10IOIIII:=IO1Il1I0OOOOIl0IOO011l1I0111OIIIII;END;PROCEDURE IIOOO0OOIll110IlI1111I1001I01IIIII(IO00lII1lIll0OllOlI1l1O0OI100IIIII:IN INTEGER;IIII1llIll1l01O1l1O0OIlO1l00OIIIII:IN INTEGER;II10ll00IlO1IIOIOIO10II0lI1l0IIIII:IN
 STD_LOGIC_VECTOR;IOIIOIIO1lIIOOl0IlO11I00II110IIIII:IN STD_LOGIC_VECTOR;II0Ol0OI111lIO001O0IIlO110IlIOIIII:OUT STD_LOGIC_VECTOR;II1ll00lO01110lOI1I0IOO0IlO0IIIIII:OUT STD_LOGIC;IO0I011OOl0OOO000O0I0O0OO0OllIIIII:OUT STD_LOGIC;IO1OllI0IIll0OIOI1l01I010OOIOOIIII:OUT
 STD_LOGIC)IS CONSTANT IIOl11l1l101llOl0l0l101I1O1llIIIII:INTEGER:=IIII1llIll1l01O1l1O0OIlO1l00OIIIII;CONSTANT III1O0Ol0IOOO0IllIOOO000O1lO0IIIII:INTEGER:=IO00lII1lIll0OllOlI1l1O0OI100IIIII-IIII1llIll1l01O1l1O0OIlO1l00OIIIII;CONSTANT IIl1IIO111llI0l1O1OI00lIl1I0OIIIII:INTEGER:=2**(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1)-1;CONSTANT IIIOOI1II1O11lOIOlOIlOOII1010IIIII:INTEGER
:=2-2**(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1);CONSTANT IO0I0I00IO00I1O0I0O0OIOOOI11IOIIII:INTEGER:=2**(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1)-1;VARIABLE IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII,IOOI0OO0l1O1O000lO10OOllOIIIIOIIII,IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:SIGNED(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+1 DOWNTO 0);VARIABLE IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII,IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII,II10110Oll1OOlIOlOlIl01111IlOIIIII:STD_LOGIC_VECTOR(IIOl11l1l101llOl0l0l101I1O1llIIIII
-1 DOWNTO 0);VARIABLE IOIO00lO11l0IOO1l0I101I11l1OOIIIII,IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII,II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII:STD_LOGIC;VARIABLE IIlO0l11I10OOIl000I0OOIO0IO0IIIIII:STD_LOGIC_VECTOR(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1 DOWNTO 0);VARIABLE IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII:STD_LOGIC_VECTOR(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1
 DOWNTO 0);VARIABLE IOIlllIIlI1OlI0l101llI0II1O1IOIIII:STD_LOGIC;VARIABLE IOO0IO0OOOOO0I10II0llO10ll1OlIIIII:STD_LOGIC_VECTOR(IIOl11l1l101llOl0l0l101I1O1llIIIII DOWNTO 0);VARIABLE IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII:STD_LOGIC_VECTOR(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+1+IIOl11l1l101llOl0l0l101I1O1llIIIII DOWNTO 0):=(
OTHERS=>'0');VARIABLE IOl10OI01O100l1IIIl0IIl1lO10lIIIII:STD_LOGIC_VECTOR(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+1+IIOl11l1l101llOl0l0l101I1O1llIIIII DOWNTO 0):=(OTHERS=>'1');VARIABLE IOI1l0OI1IO0llll1llO11Ol1IIlIIIIII:STD_LOGIC;VARIABLE IO00l1II1l000l0I11O010I1IlOlIOIIII:
STD_LOGIC;VARIABLE II0IO0O1III0I1I1OlI0011O001IOIIIII:STD_LOGIC;VARIABLE IIl1OOO111O0O11l1OOllOIIIIIl0IIIII:STD_LOGIC;VARIABLE IO00O1llIl1l1I1IIOl11OIlI1lIOOIIII:STD_LOGIC;VARIABLE IOl1I001lIl1Il1I11lI00l11O1OOIIIII:STD_LOGIC;VARIABLE
 IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII:BOOLEAN;VARIABLE III0l0O0I11OOO1lI0OOIO0llOlIlIIIII:BOOLEAN;VARIABLE IOO01101I01OlOIO111IIl0OOIOI0IIIII:BOOLEAN;VARIABLE II00l0IOI1lIlOlOOI0I011O1110OIIIII:BOOLEAN;VARIABLE IOIO1OI0IlI1I1010lO000IO01Ol0IIIII:BOOLEAN;VARIABLE IIO00Il10lI0OOllOOO0lO11lOOlIOIIII:BOOLEAN;
VARIABLE IIIIOOlIIO11011I1IlOO10OOOO0OIIIII:BOOLEAN;VARIABLE IIO0101IlI11I0IOlI01l1ll0O10OIIIII:BOOLEAN;VARIABLE IOl00OIO0IOOllO1I1O101lIIl11OIIIII:BOOLEAN;VARIABLE IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII:STD_LOGIC;VARIABLE IO00OI0ll1l1l0llI1I000OOO0010IIIII:STD_LOGIC;VARIABLE IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII
:STD_LOGIC;VARIABLE IOI0111Il0IllIIO0O0lO0I111010IIIII:STD_LOGIC;VARIABLE IOO0IOIOOll0Il0OlI001lIIIOOOIIIIII:STD_LOGIC;BEGIN IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII:=SIGNED(RESIZE(UNSIGNED(II10ll00IlO1IIOIOIO10II0lI1l0IIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO IIOl11l1l101llOl0l0l101I1O1llIIIII-1)),III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+2));IOIO00lO11l0IOO1l0I101I11l1OOIIIII:=II10ll00IlO1IIOIOIO10II0lI1l0IIIII(
IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1);IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-1 DOWNTO 0):='1'&II10ll00IlO1IIOIOIO10II0lI1l0IIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO 0);IOOI0OO0l1O1O000lO10OOllOIIIIOIIII:=SIGNED(RESIZE(UNSIGNED(IOIIOIIO1lIIOOl0IlO11I00II110IIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO IIOl11l1l101llOl0l0l101I1O1llIIIII-1)),III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+2));IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII:=IOIIOIIO1lIIOOl0IlO11I00II110IIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1);IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-1
 DOWNTO 0):='1'&IOIIOIIO1lIIOOl0IlO11I00II110IIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO 0);II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII:=(IOIO00lO11l0IOO1l0I101I11l1OOIIIII XOR IIIIl0I1lO1llIOIOOO1lOl11IIlOIIIII);IOO01101I01OlOIO111IIl0OOIOI0IIIII:=FLT_PT_IS_INF(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,II10ll00IlO1IIOIOIO10II0lI1l0IIIII);IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII:=FLT_PT_IS_NAN(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,II10ll00IlO1IIOIOIO10II0lI1l0IIIII);IOIO1OI0IlI1I1010lO000IO01Ol0IIIII:=
II1IOOO1II0l1lOl00I1O001I00O0IIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,II10ll00IlO1IIOIOIO10II0lI1l0IIIII);II00l0IOI1lIlOlOOI0I011O1110OIIIII:=FLT_PT_IS_INF(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,IOIIOIIO1lIIOOl0IlO11I00II110IIIII);III0l0O0I11OOO1lI0OOIO0llOlIlIIIII:=FLT_PT_IS_NAN(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,IOIIOIIO1lIIOOl0IlO11I00II110IIIII);IIO00Il10lI0OOllOOO0lO11lOOlIOIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII
(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,IOIIOIIO1lIIOOl0IlO11I00II110IIIII);IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII:='0';IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII:='0';IO00OI0ll1l1l0llI1I000OOO0010IIIII:='0';IIIIOOlIIO11011I1IlOO10OOOO0OIIIII:=FALSE;IIO0101IlI11I0IOlI01l1ll0O10OIIIII:=FALSE;IOl00OIO0IOOllO1I1O101lIIl11OIIIII:=FALSE;IF IOlO1OI10Il1OllOl1IIOOIO0I1lIIIIII OR III0l0O0I11OOO1lI0OOIO0llOlIlIIIII THEN IIIIOOlIIO11011I1IlOO10OOOO0OIIIII:=TRUE;ELSIF(IOO01101I01OlOIO111IIl0OOIOI0IIIII AND
 IIO00Il10lI0OOllOOO0lO11lOOlIOIIII)OR(II00l0IOI1lIlOlOOI0I011O1110OIIIII AND IOIO1OI0IlI1I1010lO000IO01Ol0IIIII)THEN IIIIOOlIIO11011I1IlOO10OOOO0OIIIII:=TRUE;IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII:='1';ELSIF IOO01101I01OlOIO111IIl0OOIOI0IIIII OR II00l0IOI1lIlOlOOI0I011O1110OIIIII THEN IIO0101IlI11I0IOlI01l1ll0O10OIIIII:=TRUE;ELSIF IOIO1OI0IlI1I1010lO000IO01Ol0IIIII OR IIO00Il10lI0OOllOOO0lO11lOOlIOIIII THEN IOl00OIO0IOOllO1I1O101lIIl11OIIIII:=TRUE;ELSE
 IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:=IIlIOIlO1lO1l1I0OOOI1O1l0O0IOIIIII+IOOI0OO0l1O1O000lO10OOllOIIIIOIIII+1-IIl1IIO111llI0l1O1OI00lIl1I0OIIIII;IIlO0l11I10OOIl000I0OOIO0IO0IIIIII:=STD_LOGIC_VECTOR(UNSIGNED(IOOll1I1OO10IlOI0lOO1lOl1O10IOIIII)*UNSIGNED(IOOIOOO1OIO1O0OIIOlOOIOlI1l1lIIIII));IF IIlO0l11I10OOIl000I0OOIO0IO0IIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1)='0'THEN IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1 DOWNTO 0):=IIlO0l11I10OOIl000I0OOIO0IO0IIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-2
 DOWNTO 0)&'0';IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:=IO1IllOO0II1ll1OII0OOO10OO0I1IIIII-1;ELSE IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII:=IIlO0l11I10OOIl000I0OOIO0IO0IIIIII;END IF;IF(IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO 0)=IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO 0))THEN IOIlllIIlI1OlI0l101llI0II1O1IOIIII:='1';ELSE IOIlllIIlI1OlI0l101llI0II1O1IOIIII:='0';END IF;IF(
IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-1)='1'AND IOIlllIIlI1OlI0l101llI0II1O1IOIIII='0')OR(IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-1)='1'AND IOIlllIIlI1OlI0l101llI0II1O1IOIIII='1'AND IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII)='1')THEN IOO0IO0OOOOO0I10II0llO10ll1OlIIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1
 DOWNTO IIOl11l1l101llOl0l0l101I1O1llIIIII)),IIOl11l1l101llOl0l0l101I1O1llIIIII+1)+1);ELSE IOO0IO0OOOOO0I10II0llO10ll1OlIIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IIOIOOI1ll1O0I1011l0O1lI0IllIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+IIOl11l1l101llOl0l0l101I1O1llIIIII-1 DOWNTO IIOl11l1l101llOl0l0l101I1O1llIIIII)),IIOl11l1l101llOl0l0l101I1O1llIIIII+1));END IF;IF IOO0IO0OOOOO0I10II0llO10ll1OlIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII)='1'THEN II10110Oll1OOlIOlOlIl01111IlOIIIII:=IOO0IO0OOOOO0I10II0llO10ll1OlIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII
 DOWNTO 1);IO1IllOO0II1ll1OII0OOO10OO0I1IIIII:=IO1IllOO0II1ll1OII0OOO10OO0I1IIIII+1;ELSE II10110Oll1OOlIOlOlIl01111IlOIIIII:=IOO0IO0OOOOO0I10II0llO10ll1OlIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-1 DOWNTO 0);END IF;IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII:='0';IO00OI0ll1l1l0llI1I000OOO0010IIIII:='0';IF IO1IllOO0II1ll1OII0OOO10OO0I1IIIII<=SIGNED(IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+1 DOWNTO 0))THEN IOl00OIO0IOOllO1I1O101lIIl11OIIIII:=TRUE;IO00OI0ll1l1l0llI1I000OOO0010IIIII
:='1';ELSIF(IO1IllOO0II1ll1OII0OOO10OO0I1IIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII+1 DOWNTO III1O0Ol0IOOO0IllIOOO000O1lO0IIIII)="01"OR(STD_LOGIC_VECTOR(IO1IllOO0II1ll1OII0OOO10OO0I1IIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1 DOWNTO 0))=NOT IIlIII1OIIl0OOl00I0IlOOI1IIlOIIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1 DOWNTO 0)))THEN IIO0101IlI11I0IOlI01l1ll0O10OIIIII:=TRUE;IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII:='1';END IF
;END IF;IF IIIIOOlIIO11011I1IlOO10OOOO0OIIIII THEN II0Ol0OI111lIO001O0IIlO110IlIOIIII:=FLT_PT_GET_QUIET_NAN(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII);ELSIF IIO0101IlI11I0IOlI01l1ll0O10OIIIII THEN II0Ol0OI111lIO001O0IIlO110IlIOIIII:=FLT_PT_GET_INF(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII);ELSIF IOl00OIO0IOOllO1I1O101lIIl11OIIIII THEN II0Ol0OI111lIO001O0IIlO110IlIOIIII:=
FLT_PT_GET_ZERO(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII,IIOl11l1l101llOl0l0l101I1O1llIIIII,II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII);ELSE II0Ol0OI111lIO001O0IIlO110IlIOIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII+III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1 DOWNTO 0):=II0l0O0IOlIOI00OIl0IlOlI01OI1IIIII&STD_LOGIC_VECTOR(IO1IllOO0II1ll1OII0OOO10OO0I1IIIII(III1O0Ol0IOOO0IllIOOO000O1lO0IIIII-1 DOWNTO 0))&II10110Oll1OOlIOlOlIl01111IlOIIIII(IIOl11l1l101llOl0l0l101I1O1llIIIII-2 DOWNTO 0);END IF;IO0I011OOl0OOO000O0I0O0OO0OllIIIII:=
IOl011Ol0O1Il1IIIIlIOlIl101IlIIIII;IO1OllI0IIll0OIOI1l01I010OOIOOIIII:=IO00OI0ll1l1l0llI1I000OOO0010IIIII;II1ll00lO01110lOI1I0IOO0IlO0IIIIII:=IOl0OIIOl0O00OO0lI0I0O1IO1OOIOIIII;END;PROCEDURE IOO0llOIlIO0110l1lOO01I00l1OIIIIII(IOIO0OOIOIOl0OIllO011O11O0OOIIIIII:IN INTEGER;IO0lI0OlO11O10O1III000O01l0l0IIIII:IN INTEGER;IIO1O00llO01OII1I11lIIO001lI0IIIII:IN BOOLEAN;IOIl1lI1IO111IO0OII101O1I0l0IOIIII:IN
 STD_LOGIC_VECTOR;IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII:IN STD_LOGIC_VECTOR;IO01O100lOO0IOOI000OO1lIOO1l0IIIII:OUT STD_LOGIC_VECTOR;IOl1100I00OlIllOI1I0III1O1l01IIIII:OUT STD_LOGIC;IO1OlIO1l10Ill0O11IO0I0ll1OlIIIIII:OUT STD_LOGIC;IIOIlOO1lI01O10O1Ol0OOI10110OIIIII:OUT
 STD_LOGIC)IS CONSTANT IO0II1lll1llOlO1lll1001O1IlOIOIIII:INTEGER:=IO0lI0OlO11O10O1III000O01l0l0IIIII;CONSTANT IOOO00lOlO0l0llI01lIlOOIIllIlIIIII:INTEGER:=IOIO0OOIOIOl0OIllO011O11O0OOIIIIII-IO0lI0OlO11O10O1III000O01l0l0IIIII;CONSTANT IIlIIII1lOllO0IlO11I1O01110IOIIIII:INTEGER:=2**(IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1)-1;CONSTANT II0I1I1l00l1O11OOIOIIllII10IlIIIII:INTEGER
:=2-2**(IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1);CONSTANT III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII:INTEGER:=2**(IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1)-1;CONSTANT III010I1Ol1OlOI0IO10O0000II11IIIII:SIGNED(IO0II1lll1llOlO1lll1001O1IlOIOIIII-1 DOWNTO 0):=(OTHERS=>'0');CONSTANT IOIlOO00I1I00lO00l0I00OlIO01IIIIII
:SIGNED(IO0II1lll1llOlO1lll1001O1IlOIOIIII DOWNTO 0):='1'&III010I1Ol1OlOI0IO10O0000II11IIIII;CONSTANT IIO111Il00001lO0l00lOOlI1IO10IIIII:SIGNED(IO0II1lll1llOlO1lll1001O1IlOIOIIII DOWNTO 0):=(OTHERS=>'0');CONSTANT II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII:SIGNED(IO0II1lll1llOlO1lll1001O1IlOIOIIII
 DOWNTO 0):=(OTHERS=>'0');CONSTANT IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII:SIGNED(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+3-1 DOWNTO 0):=IIO111Il00001lO0l00lOOlI1IO10IIIII&'1'&II10IOlI11OOI1IO1OlI0IlI0I0I1IIIII;CONSTANT IO0I10OO0llIIlII1I01OOI001IIIIIIII:SIGNED(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+2
 DOWNTO 0):=(OTHERS=>'0');VARIABLE II110IlI0l101IO1IlI1O00llI00OIIIII:STD_LOGIC_VECTOR(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1 DOWNTO 0);VARIABLE III0O000IO1IOIO10l0I00lOIII11IIIII:STD_LOGIC;VARIABLE II1llIOlOlll00O010O1lI1IOI1I1IIIII:
STD_LOGIC;VARIABLE IO1I11OIllI1III1III11OlIIlIIOIIIII:STD_LOGIC;VARIABLE IIl11lIlOO0IIII0IOlI0l1000I1IIIIII:SIGNED(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+2 DOWNTO 0);VARIABLE IOOI10l11llO01llIIllOI1IO0l1OIIIII:SIGNED(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+2 DOWNTO 0);VARIABLE IOO1IIll11IlI110IOlllI1Il1IO1IIIII
:INTEGER;VARIABLE IOO000O0Ol1OlIOOI00l11I1l1I00IIIII:INTEGER;VARIABLE IIll0O11l1O1lOl111IIOlOIl0I0OIIIII:INTEGER;VARIABLE IIOI10lI0II00O0IOOl0I10001lO1IIIII:STD_LOGIC;VARIABLE IIO1IIOOO0OO1100OO11l0OOllIIIOIIII:STD_LOGIC;VARIABLE IOO01O011lIIIlOl1O0lOIOOI110IOIIII:SIGNED
(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+2 DOWNTO 0);VARIABLE IOIOO101OO01Ol1101l1O01O1OOllIIIII:STD_LOGIC;VARIABLE IIOO0IIlO0O0I01l00I1011II0011IIIII:INTEGER;VARIABLE IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII:INTEGER;VARIABLE IIOlI0O00IO011lIIOl100O001lIOOIIII:BOOLEAN;VARIABLE
 III0IlIOll1Ill0I0I0OlIO10I1I1IIIII:BOOLEAN;VARIABLE IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII:BOOLEAN;VARIABLE II0I1O11OOll0l0I11O110OlI0lIOOIIII:BOOLEAN;VARIABLE II1lI1l0l00llI0l0l1O0OOII10I1IIIII:BOOLEAN;VARIABLE II0l10llII1lO0O1lOIlOOI10I0lIIIIII:BOOLEAN;BEGIN III0O000IO1IOIO10l0I00lOIII11IIIII:='0';
II1llIOlOlll00O010O1lI1IOI1I1IIIII:='0';IO1I11OIllI1III1III11OlIIlIIOIIIII:='0';IIOI10lI0II00O0IOOl0I10001lO1IIIII:=IOIl1lI1IO111IO0OII101O1I0l0IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1);IIO1IIOOO0OO1100OO11l0OOllIIIOIIII:=IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-1);IF IIO1O00llO01OII1I11lIIO001lI0IIIII THEN IIO1IIOOO0OO1100OO11l0OOllIIIOIIII:=NOT IIO1IIOOO0OO1100OO11l0OOllIIIOIIII;END IF;IIOlI0O00IO011lIIOl100O001lIOOIIII:=FLT_PT_IS_INF(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII
,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOIl1lI1IO111IO0OII101O1I0l0IOIIII);III0IlIOll1Ill0I0I0OlIO10I1I1IIIII:=FLT_PT_IS_NAN(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOIl1lI1IO111IO0OII101O1I0l0IOIIII);IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOIl1lI1IO111IO0OII101O1I0l0IOIIII);II0I1O11OOll0l0I11O110OlI0lIOOIIII:=FLT_PT_IS_INF(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII);II1lI1l0l00llI0l0l1O0OOII10I1IIIII:=
FLT_PT_IS_NAN(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII);II0l10llII1lO0O1lOIlOOI10I0lIIIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII);IF III0IlIOll1Ill0I0I0OlIO10I1I1IIIII OR II1lI1l0l00llI0l0l1O0OOII10I1IIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_QUIET_NAN(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII);
ELSIF IIOlI0O00IO011lIIOl100O001lIOOIIII AND II0I1O11OOll0l0I11O110OlI0lIOOIIII THEN IF IIOI10lI0II00O0IOOl0I10001lO1IIIII=IIO1IIOOO0OO1100OO11l0OOllIIIOIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_INF(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IIOI10lI0II00O0IOOl0I10001lO1IIIII);ELSE II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_QUIET_NAN(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII);
III0O000IO1IOIO10l0I00lOIII11IIIII:='1';END IF;ELSIF IIOlI0O00IO011lIIOl100O001lIOOIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_INF(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IIOI10lI0II00O0IOOl0I10001lO1IIIII);ELSIF II0I1O11OOll0l0I11O110OlI0lIOOIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_INF(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IIO1IIOOO0OO1100OO11l0OOllIIIOIIII);
ELSIF IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII AND II0l10llII1lO0O1lOIlOOI10I0lIIIIII THEN IF(IIOI10lI0II00O0IOOl0I10001lO1IIIII='1'AND IIO1IIOOO0OO1100OO11l0OOllIIIOIIII='1')THEN IOIOO101OO01Ol1101l1O01O1OOllIIIII:='1';ELSE IOIOO101OO01Ol1101l1O01O1OOllIIIII:='0';END IF;II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_ZERO(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,
IOIOO101OO01Ol1101l1O01O1OOllIIIII);ELSIF IOOllIl0I1ll0lII0IOIIO1lI10IIIIIII THEN IF IIO1IIOOO0OO1100OO11l0OOllIIIOIIII='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:='1'&IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO 0);ELSE II110IlI0l101IO1IlI1O00llI00OIIIII:='0'&IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO 0);END IF;ELSIF II0l10llII1lO0O1lOIlOOI10I0lIIIIII
 THEN IF IIOI10lI0II00O0IOOl0I10001lO1IIIII='1'THEN II110IlI0l101IO1IlI1O00llI00OIIIII:='1'&IOIl1lI1IO111IO0OII101O1I0l0IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO 0);ELSE II110IlI0l101IO1IlI1O00llI00OIIIII:='0'&IOIl1lI1IO111IO0OII101O1I0l0IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO 0);END IF;ELSE IIl11lIlOO0IIII0IOlI0l1000I1IIIIII:=(OTHERS=>'0');IIl11lIlOO0IIII0IOlI0l1000I1IIIIII(2
*IO0II1lll1llOlO1lll1001O1IlOIOIIII):='1';IIl11lIlOO0IIII0IOlI0l1000I1IIIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII-1 DOWNTO IO0II1lll1llOlO1lll1001O1IlOIOIIII+1):=SIGNED(IOIl1lI1IO111IO0OII101O1I0l0IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII-2 DOWNTO 0));IOO1IIll11IlI110IOlllI1Il1IO1IIIII:=TO_INTEGER(UNSIGNED(IOIl1lI1IO111IO0OII101O1I0l0IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO IO0II1lll1llOlO1lll1001O1IlOIOIIII-1)));IOO1IIll11IlI110IOlllI1Il1IO1IIIII:=IOO1IIll11IlI110IOlllI1Il1IO1IIIII-
IIlIIII1lOllO0IlO11I1O01110IOIIIII;IOOI10l11llO01llIIllOI1IO0l1OIIIII:=(OTHERS=>'0');IOOI10l11llO01llIIllOI1IO0l1OIIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII):='1';IOOI10l11llO01llIIllOI1IO0l1OIIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII-1 DOWNTO IO0II1lll1llOlO1lll1001O1IlOIOIIII+1):=SIGNED(IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII-2 DOWNTO 0));IOO000O0Ol1OlIOOI00l11I1l1I00IIIII:=TO_INTEGER(UNSIGNED(IOOIOOOlO000O1I0lOI1OO01l0OOlIIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII
+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII-2 DOWNTO IO0II1lll1llOlO1lll1001O1IlOIOIIII-1)));IOO000O0Ol1OlIOOI00l11I1l1I00IIIII:=IOO000O0Ol1OlIOOI00l11I1l1I00IIIII-IIlIIII1lOllO0IlO11I1O01110IOIIIII;IF IOO1IIll11IlI110IOlllI1Il1IO1IIIII>IOO000O0Ol1OlIOOI00l11I1l1I00IIIII THEN IIll0O11l1O1lOl111IIOlOIl0I0OIIIII:=IOO1IIll11IlI110IOlllI1Il1IO1IIIII-IOO000O0Ol1OlIOOI00l11I1l1I00IIIII;IIOO0IIlO0O0I01l00I1011II0011IIIII:=IOO1IIll11IlI110IOlllI1Il1IO1IIIII;IOOI10l11llO01llIIllOI1IO0l1OIIIII:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(IOOI10l11llO01llIIllOI1IO0l1OIIIII,
IIll0O11l1O1lOl111IIOlOIl0I0OIIIII);ELSE IIll0O11l1O1lOl111IIOlOIl0I0OIIIII:=IOO000O0Ol1OlIOOI00l11I1l1I00IIIII-IOO1IIll11IlI110IOlllI1Il1IO1IIIII;IIOO0IIlO0O0I01l00I1011II0011IIIII:=IOO000O0Ol1OlIOOI00l11I1l1I00IIIII;IIl11lIlOO0IIII0IOlI0l1000I1IIIIII:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(IIl11lIlOO0IIII0IOlI0l1000I1IIIIII,IIll0O11l1O1lOl111IIOlOIl0I0OIIIII);END IF;IF IIOI10lI0II00O0IOOl0I10001lO1IIIII='0'THEN IF IIO1IIOOO0OO1100OO11l0OOllIIIOIIII='0'THEN
 IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IIl11lIlOO0IIII0IOlI0l1000I1IIIIII+IOOI10l11llO01llIIllOI1IO0l1OIIIII;ELSE IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IIl11lIlOO0IIII0IOlI0l1000I1IIIIII-IOOI10l11llO01llIIllOI1IO0l1OIIIII;END IF;ELSE IF IIO1IIOOO0OO1100OO11l0OOllIIIOIIII='0'THEN IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IOOI10l11llO01llIIllOI1IO0l1OIIIII-IIl11lIlOO0IIII0IOlI0l1000I1IIIIII;ELSE IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=-(IIl11lIlOO0IIII0IOlI0l1000I1IIIIII+IOOI10l11llO01llIIllOI1IO0l1OIIIII);END
 IF;END IF;IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+2)='1'THEN IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=ABS(IOO01O011lIIIlOl1O0lOIOOI110IOIIII);IOIOO101OO01Ol1101l1O01O1OOllIIIII:='1';ELSE IOIOO101OO01Ol1101l1O01O1OOllIIIII:='0';END IF;IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+1)='1'THEN IOO01O011lIIIlOl1O0lOIOOI110IOIIII
:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(IOO01O011lIIIlOl1O0lOIOOI110IOIIII,1);IIOO0IIlO0O0I01l00I1011II0011IIIII:=IIOO0IIlO0O0I01l00I1011II0011IIIII+1;ELSE IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII:=0;WHILE IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII<2*IO0II1lll1llOlO1lll1001O1IlOIOIIII AND IOO01O011lIIIlOl1O0lOIOOI110IOIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII)='0'LOOP IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IOO01O011lIIIlOl1O0lOIOOI110IOIIII SLL 1
;IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII:=IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII+1;END LOOP;IIOO0IIlO0O0I01l00I1011II0011IIIII:=IIOO0IIlO0O0I01l00I1011II0011IIIII-IOl0lOIIO0IllIOIO1Oll0lOOOII1IIIII;END IF;IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII)='0'THEN ELSIF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII DOWNTO 0)=IOIlOO00I1I00lO00l0I00OlIO01IIIIII
 THEN IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(IO0II1lll1llOlO1lll1001O1IlOIOIIII+1)='1'THEN IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IOO01O011lIIIlOl1O0lOIOOI110IOIIII+IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII;ELSE END IF;ELSE IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=IOO01O011lIIIlOl1O0lOIOOI110IOIIII+IO1lO1OOOl00OOI0lOI1Ol1O1lI0IIIIII;END IF;IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII+1)='1'
THEN IOO01O011lIIIlOl1O0lOIOOI110IOIIII:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(IOO01O011lIIIlOl1O0lOIOOI110IOIIII,1);IIOO0IIlO0O0I01l00I1011II0011IIIII:=IIOO0IIlO0O0I01l00I1011II0011IIIII+1;END IF;IF IOO01O011lIIIlOl1O0lOIOOI110IOIIII=IO0I10OO0llIIlII1I01OOI001IIIIIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_ZERO(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,'0');ELSIF
 IIOO0IIlO0O0I01l00I1011II0011IIIII<II0I1I1l00l1O11OOIOIIllII10IlIIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_ZERO(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOIOO101OO01Ol1101l1O01O1OOllIIIII);IO1I11OIllI1III1III11OlIIlIIOIIIII:='1';ELSIF IIOO0IIlO0O0I01l00I1011II0011IIIII>III0lIIOOIOl0ll0ll0l1lO10IlIIIIIII THEN II110IlI0l101IO1IlI1O00llI00OIIIII:=FLT_PT_GET_INF
(IO0II1lll1llOlO1lll1001O1IlOIOIIII+IOOO00lOlO0l0llI01lIlOOIIllIlIIIII,IO0II1lll1llOlO1lll1001O1IlOIOIIII,IOIOO101OO01Ol1101l1O01O1OOllIIIII);II1llIOlOlll00O010O1lI1IOI1I1IIIII:='1';ELSE IIOO0IIlO0O0I01l00I1011II0011IIIII:=IIOO0IIlO0O0I01l00I1011II0011IIIII+IIlIIII1lOllO0IlO11I1O01110IOIIIII;II110IlI0l101IO1IlI1O00llI00OIIIII:=IOIOO101OO01Ol1101l1O01O1OOllIIIII&STD_LOGIC_VECTOR(TO_UNSIGNED(IIOO0IIlO0O0I01l00I1011II0011IIIII,IOOO00lOlO0l0llI01lIlOOIIllIlIIIII))&
STD_LOGIC_VECTOR(IOO01O011lIIIlOl1O0lOIOOI110IOIIII(2*IO0II1lll1llOlO1lll1001O1IlOIOIIII-1 DOWNTO IO0II1lll1llOlO1lll1001O1IlOIOIIII+1));END IF;END IF;IO01O100lOO0IOOI000OO1lIOO1l0IIIII:=II110IlI0l101IO1IlI1O00llI00OIIIII;IOl1100I00OlIllOI1I0III1O1l01IIIII:=III0O000IO1IOIO10l0I00lOIII11IIIII;IO1OlIO1l10Ill0O11IO0I0ll1OlIIIIII:=II1llIOlOlll00O010O1lI1IOI1I1IIIII;IIOIlOO1lI01O10O1Ol0OOI10110OIIIII:=IO1I11OIllI1III1III11OlIIlIIOIIIII
;END;PROCEDURE IO1I1OlOI1OII110llI1lI0IIl0O0IIIII(II110IO0lllI1lOI110IO00I1lOlIIIIII:IN INTEGER;IIl110lllO10l0llOI11l01I0I1OlIIIII:IN INTEGER;IOOll11IO1O1llOIl10010O1IIOOIIIIII:IN INTEGER;IIII00I101O111lII1O000IO1lOOIIIIII:IN INTEGER;IOOI01II11O1I1IOII1II01O1001lIIIII:IN STD_LOGIC_VECTOR;IO111Il1I1O0lO1OlOI0l01I1O010IIIII:OUT
 STD_LOGIC_VECTOR;III011IIIl1IO1l0O11000I0llI00IIIII:OUT STD_LOGIC;II1O1ll0lOO0Ol1O0OO01I0OI0lIIOIIII:OUT STD_LOGIC;IIO1l1Ol1l11Il0000II00lI011I0IIIII:OUT STD_LOGIC)IS CONSTANT IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII:INTEGER:=II110IO0lllI1lOI110IO00I1lOlIIIIII-IIl110lllO10l0llOI11l01I0I1OlIIIII;
CONSTANT II1lI11lI1II1000lOllIOl01l0l0IIIII:INTEGER:=IOOll11IO1O1llOIl10010O1IIOOIIIIII-IIII00I101O111lII1O000IO1lOOIIIIII;CONSTANT II0l0001lI0I0IlllI1I100OO10IIIIIII:INTEGER:=2**(IIO1OllIOO1lI1OOO1IOIII1lIl0IOIIII-1)-1;CONSTANT II01l0llO10l10II111lIlOIllO0lIIIII:INTEGER:=2**(II1lI11lI1II1000lOllIOl01l0l0IIIII-1)-
1;CONSTANT IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII:INTEGER:=2-2**(II1lI11lI1II1000lOllIOl01l0l0IIIII-1);CONSTANT IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII:INTEGER:=2**(II1lI11lI1II1000lOllIOl01l0l0IIIII-1)-1;CONSTANT IIl1O01ll1111l0llIOO0OOl1ll0IOIIII:UNSIGNED(
IIl110lllO10l0llOI11l01I0I1OlIIIII-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE II10l111IOllO0O1111Ill001lll1IIIII:STD_LOGIC;VARIABLE IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII:STD_LOGIC;VARIABLE IIll1lO0l0lI0OII00l00OO11IlO1IIIII:STD_LOGIC;VARIABLE
 III00O11l11IlIOI1llIIIOII100lIIIII:BOOLEAN;VARIABLE IO1l01O110OIl00l10lOOlI0lI0I0IIIII:BOOLEAN;VARIABLE IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII:BOOLEAN;VARIABLE IOIIOO1001lI01IOOlOllIOOIO1O1IIIII:UNSIGNED(IIl110lllO10l0llOI11l01I0I1OlIIIII DOWNTO 0);VARIABLE IIOlIO1l10OOO1l1IlII1ll0100IOIIIII:
INTEGER;VARIABLE III1I01Ill1l0lOIlO01lO0I1IlIIOIIII:STD_LOGIC;VARIABLE IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII:BOOLEAN;VARIABLE IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:INTEGER;VARIABLE III11I01Ol11IOO00IOI1I11OOl10IIIII:UNSIGNED(IIII00I101O111lII1O000IO1lOOIIIIII DOWNTO 0);
VARIABLE IIl1lOIllIlIl01ll00O11OIl100IOIIII:BOOLEAN:=FALSE;VARIABLE IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:STD_LOGIC_VECTOR(IOOll11IO1O1llOIl10010O1IIOOIIIIII-1 DOWNTO 0);BEGIN II10l111IOllO0O1111Ill001lll1IIIII:='0';IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII:='0';
IIll1lO0l0lI0OII00l00OO11IlO1IIIII:='0';III1I01Ill1l0lOIlO01lO0I1IlIIOIIII:=IOOI01II11O1I1IOII1II01O1001lIIIII(II110IO0lllI1lOI110IO00I1lOlIIIIII-1);III00O11l11IlIOI1llIIIOII100lIIIII:=FLT_PT_IS_INF(II110IO0lllI1lOI110IO00I1lOlIIIIII,IIl110lllO10l0llOI11l01I0I1OlIIIII,IOOI01II11O1I1IOII1II01O1001lIIIII);IO1l01O110OIl00l10lOOlI0lI0I0IIIII:=FLT_PT_IS_NAN(II110IO0lllI1lOI110IO00I1lOlIIIIII,IIl110lllO10l0llOI11l01I0I1OlIIIII,IOOI01II11O1I1IOII1II01O1001lIIIII);IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII:=
II1IOOO1II0l1lOl00I1O001I00O0IIIII(II110IO0lllI1lOI110IO00I1lOlIIIIII,IIl110lllO10l0llOI11l01I0I1OlIIIII,IOOI01II11O1I1IOII1II01O1001lIIIII);IF IO1l01O110OIl00l10lOOlI0lI0I0IIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=FLT_PT_GET_QUIET_NAN(IOOll11IO1O1llOIl10010O1IIOOIIIIII,IIII00I101O111lII1O000IO1lOOIIIIII);ELSIF III00O11l11IlIOI1llIIIOII100lIIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=
FLT_PT_GET_INF(IOOll11IO1O1llOIl10010O1IIOOIIIIII,IIII00I101O111lII1O000IO1lOOIIIIII,III1I01Ill1l0lOIlO01lO0I1IlIIOIIII);ELSIF IIlIO1lIl0lI1lOlI0I0O0I0OO0IIIIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=FLT_PT_GET_ZERO(IOOll11IO1O1llOIl10010O1IIOOIIIIII,IIII00I101O111lII1O000IO1lOOIIIIII,III1I01Ill1l0lOIlO01lO0I1IlIIOIIII);ELSIF IIII00I101O111lII1O000IO1lOOIIIIII=
IIl110lllO10l0llOI11l01I0I1OlIIIII AND IOOll11IO1O1llOIl10010O1IIOOIIIIII=II110IO0lllI1lOI110IO00I1lOlIIIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=IOOI01II11O1I1IOII1II01O1001lIIIII;ELSE IOIIOO1001lI01IOOlOllIOOIO1O1IIIII:=UNSIGNED("01"&IOOI01II11O1I1IOII1II01O1001lIIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII-2 DOWNTO 0));IIOlIO1l10OOO1l1IlII1ll0100IOIIIII:=TO_INTEGER(UNSIGNED(IOOI01II11O1I1IOII1II01O1001lIIIII(II110IO0lllI1lOI110IO00I1lOlIIIIII-2 DOWNTO IIl110lllO10l0llOI11l01I0I1OlIIIII-1
)));IIOlIO1l10OOO1l1IlII1ll0100IOIIIII:=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII-II0l0001lI0I0IlllI1I100OO10IIIIIII;IF IIl110lllO10l0llOI11l01I0I1OlIIIII<IIII00I101O111lII1O000IO1lOOIIIIII THEN III11I01Ol11IOO00IOI1I11OOl10IIIII(IIII00I101O111lII1O000IO1lOOIIIIII DOWNTO IIII00I101O111lII1O000IO1lOOIIIIII-IIl110lllO10l0llOI11l01I0I1OlIIIII):=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII DOWNTO 0);III11I01Ol11IOO00IOI1I11OOl10IIIII(IIII00I101O111lII1O000IO1lOOIIIIII
-IIl110lllO10l0llOI11l01I0I1OlIIIII-1 DOWNTO 0):=(OTHERS=>'0');IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII;ELSE IF IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII>1 THEN IIl1lOIllIlIl01ll00O11OIl100IOIIII:=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII-2 DOWNTO 0)=IIl1O01ll1111l0llIOO0OOl1ll0IOIIII(
IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII-2 DOWNTO 0);ELSE IIl1lOIllIlIl01ll00O11OIl100IOIIII:=TRUE;END IF;IF IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII>0 THEN IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII:=(IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII-1)='1')AND(NOT(IIl1lOIllIlIl01ll00O11OIl100IOIIII)OR(
IIl1lOIllIlIl01ll00O11OIl100IOIIII AND(IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII)='1')));IF IOOIl1OOO1IIl11O00lI1IlOIIl0OIIIII THEN III11I01Ol11IOO00IOI1I11OOl10IIIII:=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII DOWNTO IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII)+1;ELSE III11I01Ol11IOO00IOI1I11OOl10IIIII:=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII(IIl110lllO10l0llOI11l01I0I1OlIIIII
 DOWNTO IIl110lllO10l0llOI11l01I0I1OlIIIII-IIII00I101O111lII1O000IO1lOOIIIIII);END IF;IF III11I01Ol11IOO00IOI1I11OOl10IIIII(IIII00I101O111lII1O000IO1lOOIIIIII)='1'THEN IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII+1;ELSE IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII;END IF;ELSE IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:=IIOlIO1l10OOO1l1IlII1ll0100IOIIIII;
III11I01Ol11IOO00IOI1I11OOl10IIIII:=IOIIOO1001lI01IOOlOllIOOIO1O1IIIII;END IF;END IF;IF IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII<IOl0I1O0OllIl0lI1IlO0OIlII0lIIIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=FLT_PT_GET_ZERO(IOOll11IO1O1llOIl10010O1IIOOIIIIII,IIII00I101O111lII1O000IO1lOOIIIIII,III1I01Ill1l0lOIlO01lO0I1IlIIOIIII);IIll1lO0l0lI0OII00l00OO11IlO1IIIII:='1';ELSIF
 IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII>IIlI1l00I0IOl1l1O0llllO0I1I0IIIIII THEN IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=FLT_PT_GET_INF(IOOll11IO1O1llOIl10010O1IIOOIIIIII,IIII00I101O111lII1O000IO1lOOIIIIII,III1I01Ill1l0lOIlO01lO0I1IlIIOIIII);IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII:='1';ELSE IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII:=IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII+II01l0llO10l10II111lIlOIllO0lIIIII;IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII:=
III1I01Ill1l0lOIlO01lO0I1IlIIOIIII&STD_LOGIC_VECTOR(TO_UNSIGNED(IOlI00ll1I0I1ll0ll01l1OOl0IlIIIIII,II1lI11lI1II1000lOllIOl01l0l0IIIII))&STD_LOGIC_VECTOR(III11I01Ol11IOO00IOI1I11OOl10IIIII(IIII00I101O111lII1O000IO1lOOIIIIII-2 DOWNTO 0));END IF;END IF;IO111Il1I1O0lO1OlOI0l01I1O010IIIII:=IIOII0OO1Ol0lOOlO1O1OOlllIllOIIIII;
III011IIIl1IO1l0O11000I0llI00IIIII:=II10l111IOllO0O1111Ill001lll1IIIII;II1O1ll0lOO0Ol1O0OO01I0OI0lIIOIIII:=IIlOI1II1OOlOl00Ol01IOl0OO0OOIIIII;IIO1l1Ol1l11Il0000II00lI011I0IIIII:=IIll1lO0l0lI0OII00l00OO11IlO1IIIII;END;PROCEDURE II1011l1lI11IlIlI0l0l00100lO0IIIII(IO1OO10IOIO11O10IOOOllllI1Il0IIIII:IN INTEGER;II1IOl1011OlI0O00l1O10OlllOI0IIIII:IN INTEGER;
IO1OIOllI1llI01O00IIl0O111IIOOIIII:IN INTEGER;IO01001lO000lI1lI0IO11lO0I1OlIIIII:IN INTEGER;IOOl11OIOl101I1I1I00lIlIlO00IIIIII:IN STD_LOGIC_VECTOR;IIlOOO01III1O0O0IOII0I0lOlIlOIIIII:OUT STD_LOGIC_VECTOR;IIIl1IO0lOOOIIlOOllOl010IOl1IOIIII:OUT STD_LOGIC;IIl010l00OlI0lO1OO11Il10lIOIOOIIII:OUT
 STD_LOGIC;IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII:OUT STD_LOGIC)IS CONSTANT IIl111Il0IIlOIO000I01l00l0111IIIII:INTEGER:=2**(IO1OO10IOIO11O10IOOOllllI1Il0IIIII-II1IOl1011OlI0O00l1O10OlllOI0IIIII-1)-1;CONSTANT II1111O0III10O0OOlOlOO1l1I1l0IIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO 0):=(
OTHERS=>'0');CONSTANT III00011101l1O1OOI0l0Il0l1l10IIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO 0):=(OTHERS=>'1');CONSTANT IO0lll11llOIOOIOI1lOOIOl000I0IIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO 0):='1'&II1111O0III10O0OOlOlOO1l1I1l0IIIII
(IO1OIOllI1llI01O00IIl0O111IIOOIIII-2 DOWNTO 0);CONSTANT IO00OO00lIlIO00llOIll10l0ll1OIIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO 0):='0'&III00011101l1O1OOI0l0Il0l1l10IIIII(IO1OIOllI1llI01O00IIl0O111IIOOIIII-2 DOWNTO 0);CONSTANT IIO1lO000Il1O0lOII1IO0OOOIO00IIIII:SIGNED
(II1IOl1011OlI0O00l1O10OlllOI0IIIII-1 DOWNTO 0):=(OTHERS=>'0');CONSTANT II1001l0I11O0IIOIl01I1ll0O0OlIIIII:SIGNED(II1IOl1011OlI0O00l1O10OlllOI0IIIII DOWNTO 0):='1'&IIO1lO000Il1O0lOII1IO0OOOIO00IIIII;CONSTANT II1II1OO1ll10IlO0I10O0OI000IIOIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII
 DOWNTO 0):=(OTHERS=>'0');CONSTANT IOOl01OO110II1I0lIlI001II11I0IIIII:SIGNED(II1IOl1011OlI0O00l1O10OlllOI0IIIII-1 DOWNTO 0):=(OTHERS=>'0');CONSTANT II0IIlIOII0IIl1lIO1llO1O1lOlIIIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII+II1IOl1011OlI0O00l1O10OlllOI0IIIII+1
 DOWNTO 0):=II1II1OO1ll10IlO0I10O0OI000IIOIIII&'1'&IOOl01OO110II1I0lIlI001II11I0IIIII;VARIABLE IIll0I0ll1ll1O0IOlO1O01llII00IIIII:SIGNED(IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO 0);VARIABLE II1ll1Il1Il11O10OllIl0l1l1l0IOIIII:STD_LOGIC;VARIABLE III0II00l1IIlIO100l00OlI1l1O0IIIII
:STD_LOGIC;VARIABLE II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:SIGNED(II1IOl1011OlI0O00l1O10OlllOI0IIIII+IO1OIOllI1llI01O00IIl0O111IIOOIIII+1 DOWNTO 0);VARIABLE IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII:INTEGER;VARIABLE III101l00lllOOOlIO0OO1lI1OO1OIIIII:INTEGER;VARIABLE II0l0l0II0Il010II1l000011O1lIIIIII:STD_LOGIC
;VARIABLE IIlIIOOI1lOO0O0I1O1O10lI0OlIOOIIII:INTEGER;CONSTANT IOO0lOOOll1OI0OI0lI10IOOOII00IIIII:SIGNED(II1IOl1011OlI0O00l1O10OlllOI0IIIII-1 DOWNTO 0):=(OTHERS=>'0');BEGIN II1ll1Il1Il11O10OllIl0l1l1l0IOIIII:='0';III0II00l1IIlIO100l00OlI1l1O0IIIII:='0';II0l0l0II0Il010II1l000011O1lIIIIII:=IOOl11OIOl101I1I1I00lIlIlO00IIIIII(
IO1OO10IOIO11O10IOOOllllI1Il0IIIII-1);IF II1IOOO1II0l1lOl00I1O001I00O0IIIII(IO1OO10IOIO11O10IOOOllllI1Il0IIIII,II1IOl1011OlI0O00l1O10OlllOI0IIIII,IOOl11OIOl101I1I1I00lIlIlO00IIIIII)THEN IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=II1111O0III10O0OOlOlOO1l1I1l0IIIII;ELSIF FLT_PT_IS_NAN(IO1OO10IOIO11O10IOOOllllI1Il0IIIII,II1IOl1011OlI0O00l1O10OlllOI0IIIII,IOOl11OIOl101I1I1I00lIlIlO00IIIIII)THEN IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=IO0lll11llOIOOIOI1lOOIOl000I0IIIII;II1ll1Il1Il11O10OllIl0l1l1l0IOIIII
:='1';ELSIF FLT_PT_IS_INF(IO1OO10IOIO11O10IOOOllllI1Il0IIIII,II1IOl1011OlI0O00l1O10OlllOI0IIIII,IOOl11OIOl101I1I1I00lIlIlO00IIIIII)THEN IF II0l0l0II0Il010II1l000011O1lIIIIII='0'THEN IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=IO00OO00lIlIO00llOIll10l0ll1OIIIII;ELSE IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=IO0lll11llOIOOIOI1lOOIOl000I0IIIII;END IF;III0II00l1IIlIO100l00OlI1l1O0IIIII:='1';II1ll1Il1Il11O10OllIl0l1l1l0IOIIII
:='1';ELSE II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:=(OTHERS=>'0');II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+IO1OIOllI1llI01O00IIl0O111IIOOIIII):='1';II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO IO1OIOllI1llI01O00IIl0O111IIOOIIII+1):=SIGNED(IOOl11OIOl101I1I1I00lIlIlO00IIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII-2 DOWNTO 0));IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII
:=TO_INTEGER(UNSIGNED(IOOl11OIOl101I1I1I00lIlIlO00IIIIII(IO1OO10IOIO11O10IOOOllllI1Il0IIIII-2 DOWNTO II1IOl1011OlI0O00l1O10OlllOI0IIIII-1)));IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII:=IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII-IIl111Il0IIlOIO000I01l00l0111IIIII;III101l00lllOOOlIO0OO1lI1OO1OIIIII:=(IO1OIOllI1llI01O00IIl0O111IIOOIIII-(IO01001lO000lI1lI0IO11lO0I1OlIIIII+1))-IOl0lI0l0O1IlOIlI1IlO1l01Il00IIIII;IF III101l00lllOOOlIO0OO1lI1OO1OIIIII>0 OR(
III101l00lllOOOlIO0OO1lI1OO1OIIIII=0 AND II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+IO1OIOllI1llI01O00IIl0O111IIOOIIII-1 DOWNTO II1IOl1011OlI0O00l1O10OlllOI0IIIII+1)=IOO0lOOOll1OI0OI0lI10IOOOII00IIIII)THEN II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(II11OIIIO0I0OI0IIIIO1lOO011IlIIIII,III101l00lllOOOlIO0OO1lI1OO1OIIIII);ELSE III0II00l1IIlIO100l00OlI1l1O0IIIII:='1';END IF;IF(
II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII)='0')THEN ELSIF II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII DOWNTO 0)=II1001l0I11O0IIOIl01I1ll0O0OlIIIII THEN IF(II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+1)='1')THEN II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:=II11OIIIO0I0OI0IIIIO1lOO011IlIIIII+II0IIlIOII0IIl1lIO1llO1O1lOlIIIIII;ELSE END IF;ELSE
 II11OIIIO0I0OI0IIIIO1lOO011IlIIIII:=II11OIIIO0I0OI0IIIIO1lOO011IlIIIII+II0IIlIOII0IIl1lIO1llO1O1lOlIIIIII;END IF;IF II0l0l0II0Il010II1l000011O1lIIIIII='1'THEN II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(IO1OIOllI1llI01O00IIl0O111IIOOIIII+II1IOl1011OlI0O00l1O10OlllOI0IIIII+1 DOWNTO II1IOl1011OlI0O00l1O10OlllOI0IIIII+1):=-II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(IO1OIOllI1llI01O00IIl0O111IIOOIIII+II1IOl1011OlI0O00l1O10OlllOI0IIIII+1 DOWNTO II1IOl1011OlI0O00l1O10OlllOI0IIIII+1);END IF;IF
(II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+1+IO1OIOllI1llI01O00IIl0O111IIOOIIII)XOR II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(II1IOl1011OlI0O00l1O10OlllOI0IIIII+IO1OIOllI1llI01O00IIl0O111IIOOIIII))='1'THEN III0II00l1IIlIO100l00OlI1l1O0IIIII:='1';END IF;IF II1ll1Il1Il11O10OllIl0l1l1l0IOIIII='1'OR III0II00l1IIlIO100l00OlI1l1O0IIIII='1'THEN IF II0l0l0II0Il010II1l000011O1lIIIIII='0'THEN
 IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=IO00OO00lIlIO00llOIll10l0ll1OIIIII;ELSE IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=IO0lll11llOIOOIOI1lOOIOl000I0IIIII;END IF;ELSE IIll0I0ll1ll1O0IOlO1O01llII00IIIII:=II11OIIIO0I0OI0IIIIO1lOO011IlIIIII(IO1OIOllI1llI01O00IIl0O111IIOOIIII+II1IOl1011OlI0O00l1O10OlllOI0IIIII DOWNTO II1IOl1011OlI0O00l1O10OlllOI0IIIII+1);END IF;END IF;IIlOOO01III1O0O0IOII0I0lOlIlOIIIII:=STD_LOGIC_VECTOR
(IIll0I0ll1ll1O0IOlO1O01llII00IIIII);IIIl1IO0lOOOIIlOOllOl010IOl1IOIIII:=II1ll1Il1Il11O10OllIl0l1l1l0IOIIII;IIl010l00OlI0lO1OO11Il10lIOIOOIIII:=III0II00l1IIlIO100l00OlI1l1O0IIIII;IIOIl1I10OOOllIlIOl11lI0IO1lIOIIII:='0';END;PROCEDURE II111O1llOOlI0lOOIIIl0OIlIlllIIIII(IIO11lIl110IO0lO00IOOl0Il11I1IIIII:IN INTEGER;II1IO0OO0IOlO11110OOlO1O0101IOIIII:IN INTEGER;
II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII:IN INTEGER;IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII:IN INTEGER;IO0lllOII000O01100OOI0II1II01IIIII:IN STD_LOGIC_VECTOR;IO0IllIIO11IlI1010IIl0l000001IIIII:OUT STD_LOGIC_VECTOR;II1l0I0l10l0I1I1lO01l10I01lI1IIIII:OUT STD_LOGIC;IIO001lIl0II1lI10I1000O00Ol10IIIII:OUT
 STD_LOGIC;IIOI1lO0I00III00II0IO0ll0111IOIIII:OUT STD_LOGIC)IS CONSTANT III11OII1IlIl1001I1IO1111l0IlIIIII:INTEGER:=II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII-IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII;CONSTANT IIII11lI1lOl0OlOO0II11lI101lOIIIII:INTEGER:=2**(III11OII1IlIl1001I1IO1111l0IlIIIII-1)-1;CONSTANT
 IOl0Ill1OOl0O1IO1l0010I0lO010IIIII:INTEGER:=0;CONSTANT IO0IlOI1OIOO0l101l10IO00l0101IIIII:INTEGER:=2**III11OII1IlIl1001I1IO1111l0IlIIIII-1;CONSTANT IIOO1OlIO01I00l0OO0I11OII1OlOIIIII:INTEGER:=FLT_PT_MAX(IIO11lIl110IO0lO00IOOl0Il11I1IIIII+1,IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII+1);CONSTANT IIOOI1O1lllllI10ll0I0OIO1IIlIIIIII:
SIGNED(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII:INTEGER;VARIABLE IIl1O1IllII0I01IlO01l0lII0lIOOIIII:SIGNED(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1 DOWNTO 0);VARIABLE IOI1IOl0OI0O1OllO10lO1lOOl0l1IIIII:
STD_LOGIC_VECTOR(II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII-1 DOWNTO 0);VARIABLE IIII00IOl0llO0O011llO1lOOOIIOIIIII:SIGNED(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1 DOWNTO 0);VARIABLE IIlOIl110lOl10lO1OIllII10IOO1IIIII:INTEGER;VARIABLE IO0O00IOlOOIOO11lI01l000IIIIOIIIII:STD_LOGIC;
VARIABLE II10I1011llOIIlI00OI0IIIl0OIOIIIII:INTEGER;VARIABLE IOI0O1l0101lI100OIOIlll001OO1IIIII:BOOLEAN;BEGIN IO0O00IOlOOIOO11lI01l000IIIIOIIIII:=IO0lllOII000O01100OOI0II1II01IIIII(IIO11lIl110IO0lO00IOOl0Il11I1IIIII-1);IIII00IOl0llO0O011llO1lOOOIIOIIIII:=(OTHERS=>'0');IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1 DOWNTO IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-IIO11lIl110IO0lO00IOOl0Il11I1IIIII-1):=
RESIZE(SIGNED(IO0lllOII000O01100OOI0II1II01IIIII),IIO11lIl110IO0lO00IOOl0Il11I1IIIII+1);IF IIOO1OlIO01I00l0OO0I11OII1OlOIIIII>(IIO11lIl110IO0lO00IOOl0Il11I1IIIII+1)THEN IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-IIO11lIl110IO0lO00IOOl0Il11I1IIIII-2 DOWNTO 0):=(OTHERS=>'0');END IF;IIlOIl110lOl10lO1OIllII10IOO1IIIII:=(IIO11lIl110IO0lO00IOOl0Il11I1IIIII-II1IO0OO0IOlO11110OOlO1O0101IOIIII)-1+IIII11lI1lOl0OlOO0II11lI101lOIIIII;IF
 IO0O00IOlOOIOO11lI01l000IIIIOIIIII='1'THEN IIII00IOl0llO0O011llO1lOOOIIOIIIII:=-IIII00IOl0llO0O011llO1lOOOIIOIIIII;END IF;II10I1011llOIIlI00OI0IIIl0OIOIIIII:=0;WHILE II10I1011llOIIlI00OI0IIIl0OIOIIIII<IIOO1OlIO01I00l0OO0I11OII1OlOIIIII AND IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-2)='0'LOOP IIII00IOl0llO0O011llO1lOOOIIOIIIII:=IIII00IOl0llO0O011llO1lOOOIIOIIIII SLL 1;II10I1011llOIIlI00OI0IIIl0OIOIIIII:=
II10I1011llOIIlI00OI0IIIl0OIOIIIII+1;END LOOP;IIlOIl110lOl10lO1OIllII10IOO1IIIII:=IIlOIl110lOl10lO1OIllII10IOO1IIIII-II10I1011llOIIlI00OI0IIIl0OIOIIIII;IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII:=IIO11lIl110IO0lO00IOOl0Il11I1IIIII-IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII;IF(IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII>0)THEN IIl1O1IllII0I01IlO01l0lII0lIOOIIII:=(OTHERS=>'0');IIl1O1IllII0I01IlO01l0lII0lIOOIIII(IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII-1):=
'1';IF IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII-1)='0'THEN ELSE IOI0O1l0101lI100OIOIlll001OO1IIIII:=TRUE;IF IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII>1 THEN FOR IIlI1lIIIOI0l01l01OOII00I0O0lIIIII IN 0 TO IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII-2 LOOP IF IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIlI1lIIIOI0l01l01OOII00I0O0lIIIII)='1'THEN IOI0O1l0101lI100OIOIlll001OO1IIIII:=FALSE;END IF;
END LOOP;END IF;IF IOI0O1l0101lI100OIOIlll001OO1IIIII THEN IF IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIIIOI0l0OOO1O1ll0OOI00lI0l1IOIIII)='1'THEN IIII00IOl0llO0O011llO1lOOOIIOIIIII:=IIII00IOl0llO0O011llO1lOOOIIOIIIII+IIl1O1IllII0I01IlO01l0lII0lIOOIIII;END IF;ELSE IIII00IOl0llO0O011llO1lOOOIIOIIIII:=IIII00IOl0llO0O011llO1lOOOIIOIIIII+IIl1O1IllII0I01IlO01l0lII0lIOOIIII;END IF;END IF;IF(
IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1))='1'THEN IIII00IOl0llO0O011llO1lOOOIIOIIIII:=II1001IO0010Oll1I01lOI0I0IlIOIIIII(IIII00IOl0llO0O011llO1lOOOIIOIIIII,1);IIlOIl110lOl10lO1OIllII10IOO1IIIII:=IIlOIl110lOl10lO1OIllII10IOO1IIIII+1;END IF;END IF;ASSERT IIlOIl110lOl10lO1OIllII10IOO1IIIII>=IOl0Ill1OOl0O1IO1l0010I0lO010IIIII REPORT
"ERROR: flt_pt_fix_to_flt: Internal error, exponent is less than minimum permitted.  Please file a Xilinx Support request quoting this error message."
SEVERITY FAILURE;ASSERT IIlOIl110lOl10lO1OIllII10IOO1IIIII<=IO0IlOI1OIOO0l101l10IO00l0101IIIII REPORT
"ERROR: flt_pt_fix_to_flt: Internal error, exponent is greater than maximum permitted.  Please file a Xilinx Support request quoting this error message."
SEVERITY FAILURE;IF IIII00IOl0llO0O011llO1lOOOIIOIIIII=IIOOI1O1lllllI10ll0I0OIO1IIlIIIIII THEN IOI1IOl0OI0O1OllO10lO1lOOl0l1IIIII:=FLT_PT_GET_ZERO(II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII,IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII,'0');ELSE IIlOIl110lOl10lO1OIllII10IOO1IIIII:=IIlOIl110lOl10lO1OIllII10IOO1IIIII;IOI1IOl0OI0O1OllO10lO1lOOl0l1IIIII:=IO0O00IOlOOIOO11lI01l000IIIIOIIIII&
STD_LOGIC_VECTOR(TO_UNSIGNED(IIlOIl110lOl10lO1OIllII10IOO1IIIII,II0lIlIIOl0I0Ol0lIl0111l1I1l1IIIII-IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII))&STD_LOGIC_VECTOR(IIII00IOl0llO0O011llO1lOOOIIOIIIII(IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-3 DOWNTO IIOO1OlIO01I00l0OO0I11OII1OlOIIIII-1-IO0OIl1OO10lO00IlIl0Il0l1l1OIIIIII));END IF;IO0IllIIO11IlI1010IIl0l000001IIIII:=IOI1IOl0OI0O1OllO10lO1lOOl0l1IIIII;
II1l0I0l10l0I1I1lO01l10I01lI1IIIII:='0';IIO001lIl0II1lI10I1000O00Ol10IIIII:='0';IIOI1lO0I00III00II0IO0ll0111IOIIII:='0';END;PROCEDURE IO1lII1OIl0llIl0IIlIlOI10l0OlIIIII(IIl000O0IO0llO0II1lI1010lOO0IOIIII:IN INTEGER;IOlO1l1O00OIII1I0l0lOll0IOlO0IIIII:IN INTEGER;IOlIll0lIIOlIl1l1lI01OII11lOIIIIII:IN INTEGER;II1OO01O01O10l0IIOIII101O1000IIIII
:IN STD_LOGIC_VECTOR(FLT_PT_COMPARE_OPERATION_WIDTH-1 DOWNTO 0);II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII:IN STD_LOGIC_VECTOR;II0I00l0IOOO11I1l0O11O1I1O101IIIII:IN STD_LOGIC_VECTOR;IOlO0lIIlI010OIO10l11l1l1lIO0IIIII:OUT STD_LOGIC_VECTOR;
II10010II0ll0l10O0OOI01I11110IIIII:OUT STD_LOGIC)IS CONSTANT IIllIl0lIO10011Ol0O10l01O1Il0IIIII:INTEGER:=IOlO1l1O00OIII1I0l0lOll0IOlO0IIIII;CONSTANT III0lIIl1lO0OI1OlO101lI10lIIIOIIII:INTEGER:=IIl000O0IO0llO0II1lI1010lOO0IOIIII-IOlO1l1O00OIII1I0l0lOll0IOlO0IIIII;CONSTANT IIO01II0O1OlI01l11l10Il10llI0IIIII:INTEGER:=2**(III0lIIl1lO0OI1OlO101lI10lIIIOIIII-1)-1;VARIABLE
 IIII10l0Ol001IlOlO1OO1l1llO00IIIII:UNSIGNED(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0);VARIABLE IO11OI1l0l1I1IOl1Ol0lIlIlOlO1IIIII:UNSIGNED(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0);VARIABLE II0lIllO11Ill0l10OIOI01I00I1OIIIII:UNSIGNED(III0lIIl1lO0OI1OlO101lI10lIIIOIIII-1 DOWNTO 0);VARIABLE IOO11lOOlO1lO1OOIIIOOl0l00OOIOIIII:UNSIGNED
(III0lIIl1lO0OI1OlO101lI10lIIIOIIII-1 DOWNTO 0);VARIABLE IOI1I0l0OllIO01I0O1O001I0lI1IOIIII:STD_LOGIC;VARIABLE II1I01lOI10OOOlO0lO1O0OOIOlI0IIIII:STD_LOGIC;VARIABLE IIIO01IOl00Il00111I010ll11010IIIII:BOOLEAN;VARIABLE IO000l1I110IOlI1l1OlO00l1011IIIIII:BOOLEAN;VARIABLE II1l1I00I1OI1Il0l111OOI10l1lIOIIII:
BOOLEAN;VARIABLE II01Il0I0I011lOlIO11Il1l11IOlIIIII:BOOLEAN;VARIABLE IO1O0O0O00O0I0100lIl10OOIlO0OIIIII:STD_LOGIC_VECTOR(3 DOWNTO 0);VARIABLE IIlOlIIOllO0I11I1OlOIlIl1IlOOIIIII:BOOLEAN;VARIABLE IIl111OlOO0lll00IOO01OOIl1l1IIIIII:
BOOLEAN;VARIABLE IIO101OI0lOlOI1IIOllllI10O1lIIIIII:STD_LOGIC;VARIABLE IIOO0lIlIOlI0Ol010ll0lIl100IIIIIII:BOOLEAN;VARIABLE II00lO01O111Ol1OOIllOOl110OOIIIIII:BOOLEAN;VARIABLE IIO00IlOO0lO0l1OO0l00lOOI0lO0IIIII:BOOLEAN;VARIABLE III110I0l00l0lOl000OOI0I1IOlIOIIII:BOOLEAN;
VARIABLE IIOI0III1IIlI00OOOI1I100OOIIOOIIII:BOOLEAN;VARIABLE IIIIOO0llOIll1IO0lIlO0l111O0IOIIII:BOOLEAN;BEGIN IIOO0lIlIOlI0Ol010ll0lIl100IIIIIII:=FLT_PT_IS_INF(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII);II00lO01O111Ol1OOIllOOl110OOIIIIII:=FLT_PT_IS_NAN(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII);IIO00IlOO0lO0l1OO0l00lOOI0lO0IIIII:=
II1IOOO1II0l1lOl00I1O001I00O0IIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII);III110I0l00l0lOl000OOI0I1IOlIOIIII:=FLT_PT_IS_INF(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II0I00l0IOOO11I1l0O11O1I1O101IIIII);IIOI0III1IIlI00OOOI1I100OOIIOOIIII:=FLT_PT_IS_NAN(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II0I00l0IOOO11I1l0O11O1I1O101IIIII);IIIIOO0llOIll1IO0lIlO0l111O0IOIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII
(IIllIl0lIO10011Ol0O10l01O1Il0IIIII+III0lIIl1lO0OI1OlO101lI10lIIIOIIII,IIllIl0lIO10011Ol0O10l01O1Il0IIIII,II0I00l0IOOO11I1l0O11O1I1O101IIIII);IOI1I0l0OllIO01I0O1O001I0lI1IOIIII:=II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII(III0lIIl1lO0OI1OlO101lI10lIIIOIIII+IIllIl0lIO10011Ol0O10l01O1Il0IIIII-1);II0lIllO11Ill0l10OIOI01I00I1OIIIII:=UNSIGNED(II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII(III0lIIl1lO0OI1OlO101lI10lIIIOIIII+IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO IIllIl0lIO10011Ol0O10l01O1Il0IIIII-1));IF IIO00IlOO0lO0l1OO0l00lOOI0lO0IIIII THEN IIII10l0Ol001IlOlO1OO1l1llO00IIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0):=(OTHERS=>'0');ELSE IIII10l0Ol001IlOlO1OO1l1llO00IIIII
(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0):=UNSIGNED(II1l10I1lIlOIIl1lO0IO0I1OOIIlIIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0));END IF;II1I01lOI10OOOlO0lO1O0OOIOlI0IIIII:=II0I00l0IOOO11I1l0O11O1I1O101IIIII(III0lIIl1lO0OI1OlO101lI10lIIIOIIII+IIllIl0lIO10011Ol0O10l01O1Il0IIIII-1);IOO11lOOlO1lO1OOIIIOOl0l00OOIOIIII:=UNSIGNED(II0I00l0IOOO11I1l0O11O1I1O101IIIII(III0lIIl1lO0OI1OlO101lI10lIIIOIIII+IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO IIllIl0lIO10011Ol0O10l01O1Il0IIIII-1));IF IIIIOO0llOIll1IO0lIlO0l111O0IOIIII THEN IO11OI1l0l1I1IOl1Ol0lIlIlOlO1IIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII
-2 DOWNTO 0):=(OTHERS=>'0');ELSE IO11OI1l0l1I1IOl1Ol0lIlIlOlO1IIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0):=UNSIGNED(II0I00l0IOOO11I1l0O11O1I1O101IIIII(IIllIl0lIO10011Ol0O10l01O1Il0IIIII-2 DOWNTO 0));END IF;IIIO01IOl00Il00111I010ll11010IIIII:=FALSE;IO000l1I110IOlI1l1OlO00l1011IIIIII:=FALSE;II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=FALSE;
II01Il0I0I011lOlIO11Il1l11IOlIIIII:=FALSE;IIO101OI0lOlOI1IIOllllI10O1lIIIIII:='0';IF(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='0'AND II1I01lOI10OOOlO0lO1O0OOIOlI0IIIII='1')THEN II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=TRUE;ELSIF(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='1'AND II1I01lOI10OOOlO0lO1O0OOIOlI0IIIII='0')THEN IO000l1I110IOlI1l1OlO00l1011IIIIII:=TRUE;ELSIF(II0lIllO11Ill0l10OIOI01I00I1OIIIII
/=IOO11lOOlO1lO1OOIIIOOl0l00OOIOIIII)THEN IF(IOO11lOOlO1lO1OOIIIOOl0l00OOIOIIII>II0lIllO11Ill0l10OIOI01I00I1OIIIII)THEN IO000l1I110IOlI1l1OlO00l1011IIIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='0');II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='1');ELSE IO000l1I110IOlI1l1OlO00l1011IIIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='1');II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='0');END IF;ELSE IF
(IO11OI1l0l1I1IOl1Ol0lIlIlOlO1IIIII>IIII10l0Ol001IlOlO1OO1l1llO00IIIII)THEN IO000l1I110IOlI1l1OlO00l1011IIIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='0');II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='1');ELSE IF(IO11OI1l0l1I1IOl1Ol0lIlIlOlO1IIIII/=IIII10l0Ol001IlOlO1OO1l1llO00IIIII)THEN IO000l1I110IOlI1l1OlO00l1011IIIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='1');II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=(IOI1I0l0OllIO01I0O1O001I0lI1IOIIII='0');ELSE
 IIIO01IOl00Il00111I010ll11010IIIII:=TRUE;END IF;END IF;END IF;IF IIO00IlOO0lO0l1OO0l00lOOI0lO0IIIII AND IIIIOO0llOIll1IO0lIlO0l111O0IOIIII THEN IIIO01IOl00Il00111I010ll11010IIIII:=TRUE;IO000l1I110IOlI1l1OlO00l1011IIIIII:=FALSE;II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=FALSE;END IF;IF II00lO01O111Ol1OOIllOOl110OOIIIIII OR IIOI0III1IIlI00OOOI1I100OOIIOOIIII THEN
 IIIO01IOl00Il00111I010ll11010IIIII:=FALSE;IO000l1I110IOlI1l1OlO00l1011IIIIII:=FALSE;II1l1I00I1OI1Il0l111OOI10l1lIOIIII:=FALSE;II01Il0I0I011lOlIO11Il1l11IOlIIIII:=TRUE;END IF;IO1O0O0O00O0I0100lIl10OOIlO0OIIIII:=(OTHERS=>'0');IF II1OO01O01O10l0IIOIII101O1000IIIII="111"THEN IF IIIO01IOl00Il00111I010ll11010IIIII THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(0):=
'1';END IF;IF IO000l1I110IOlI1l1OlO00l1011IIIIII THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(1):='1';END IF;IF II1l1I00I1OI1Il0l111OOI10l1lIOIIII THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(2):='1';END IF;IF II01Il0I0I011lOlIO11Il1l11IOlIIIII THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(3):='1';END IF;ELSIF((
II1l1I00I1OI1Il0l111OOI10l1lIOIIII AND(II1OO01O01O10l0IIOIII101O1000IIIII(2)='1'))OR(IIIO01IOl00Il00111I010ll11010IIIII AND(II1OO01O01O10l0IIOIII101O1000IIIII(1)='1'))OR(IO000l1I110IOlI1l1OlO00l1011IIIIII AND(II1OO01O01O10l0IIOIII101O1000IIIII(0)='1')))THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(0):='1';ELSIF(II1OO01O01O10l0IIOIII101O1000IIIII="000")THEN IF
(II01Il0I0I011lOlIO11Il1l11IOlIIIII)THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(0):='1';END IF;END IF;IF(II1OO01O01O10l0IIOIII101O1000IIIII/="111"AND((II01Il0I0I011lOlIO11Il1l11IOlIIIII AND NOT(II1OO01O01O10l0IIOIII101O1000IIIII="000"OR II1OO01O01O10l0IIOIII101O1000IIIII="010"OR II1OO01O01O10l0IIOIII101O1000IIIII="101"))))THEN
 IIO101OI0lOlOI1IIOllllI10O1lIIIIII:='1';IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(0):='0';END IF;IF(II01Il0I0I011lOlIO11Il1l11IOlIIIII AND II1OO01O01O10l0IIOIII101O1000IIIII="101")THEN IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(0):='1';END IF;IF IOlIll0lIIOlIl1l1lI01OII11lOIIIIII>4 THEN IOlO0lIIlI010OIO10l11l1l1lIO0IIIII(3 DOWNTO 0):=IO1O0O0O00O0I0100lIl10OOIlO0OIIIII
;FOR IO0O1OIIlI0I0101llOI1O01OOIIOOIIII IN 4 TO IOlIll0lIIOlIl1l1lI01OII11lOIIIIII-1 LOOP IOlO0lIIlI010OIO10l11l1l1lIO0IIIII(IO0O1OIIlI0I0101llOI1O01OOIIOOIIII):='0';END LOOP;ELSE IOlO0lIIlI010OIO10l11l1l1lIO0IIIII:=IO1O0O0O00O0I0100lIl10OOIlO0OIIIII(IOlIll0lIIOlIl1l1lI01OII11lOIIIIII-1 DOWNTO 0);END IF;II10010II0ll0l10O0OOI01I11110IIIII:=IIO101OI0lOlOI1IIOllllI10O1lIIIIII;END;PROCEDURE
 IOOOOI1lIlOlI10IOOOI00O10O00IIIIII(II1O1lIOOI00OOI10010I1010IOOOIIIII:IN INTEGER;IOO0IlOlIOOll110I1l0O0011lllIOIIII:IN INTEGER;IOOl1IIO0I01ll0O00O01O1I000IOIIIII:IN STD_LOGIC_VECTOR;IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:OUT STD_LOGIC_VECTOR;III1lI0IOlOO11l0lO0IIl00OlOl0IIIII:OUT STD_LOGIC;IIO1lIlIlIIll0011II00OlO00llOIIIII:OUT
 STD_LOGIC)IS CONSTANT IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII:INTEGER:=IOO0IlOlIOOll110I1l0O0011lllIOIIII;CONSTANT IIOl00111100II1IOl0O1OO1I0lIOOIIII:INTEGER:=II1O1lIOOI00OOI10010I1010IOOOIIIII-IOO0IlOlIOOll110I1l0O0011lllIOIIII;VARIABLE II101I1OIIl111101l00ll0Ol1l01IIIII:STD_LOGIC_VECTOR(IIOl00111100II1IOl0O1OO1I0lIOOIIII-1 DOWNTO 0);VARIABLE IO1ll0OlO000O0lIO01I1llIOlOI1IIIII:
STD_LOGIC_VECTOR(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-2 DOWNTO 0);VARIABLE IOI111lOI111OOlI0III1I0lO1I0IIIIII:STD_LOGIC;VARIABLE IOl0l0l0I0I0l0I010011l0llIl1lIIIII:BOOLEAN;VARIABLE IO1l0OlOOl00O1OIlI0O0lIIlIlOlIIIII:BOOLEAN;VARIABLE II001lI100O0O0I1l1IIOlIlO00IlIIIII:BOOLEAN;VARIABLE
 IO1Ol0OlIIO11llOOl00IIIO11101IIIII:STD_LOGIC_VECTOR(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII-1 DOWNTO 0);VARIABLE IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:STD_LOGIC;VARIABLE II0O01100OIIIl10O1OIl0I00Ol10IIIII:STD_LOGIC;CONSTANT II1I1IOl0I0I1I0lIl00ll11I111OIIIII:INTEGER:=
FLT_PT_RECIP_W(IOO0IlOlIOOll110I1l0O0011lllIOIIII);CONSTANT IO0O010II00IOl10I10O1l0I10O1IOIIII:INTEGER:=FLT_PT_RECIP_K(II1O1lIOOI00OOI10010I1010IOOOIIIII,IOO0IlOlIOOll110I1l0O0011lllIOIIII,FLT_PT_RECIP_OP_CODE);CONSTANT II11OlI0I00OIO1llOI00O0lI0OlIIIIII:INTEGER:=FLT_PT_RECIP_M(II1O1lIOOI00OOI10010I1010IOOOIIIII,IOO0IlOlIOOll110I1l0O0011lllIOIIII);
CONSTANT IO1I1OO00O1lIOOIll0lIO0l10lIlIIIII:INTEGER:=(2*II11OlI0I00OIO1llOI00O0lI0OlIIIIII)+3;VARIABLE IOOlII11IOO011lOll1IOO10O010OIIIII:STD_LOGIC_VECTOR(IO0O010II00IOl10I10O1l0I10O1IOIIII-1 DOWNTO 0);VARIABLE IOI1IlOO001111I101I1O01l01lI1IIIII:STD_LOGIC_VECTOR(II11OlI0I00OIO1llOI00O0lI0OlIIIIII-1 DOWNTO
 0);VARIABLE II1l0l1O010I00O1Ill1O10lIII0OIIIII:STD_LOGIC_VECTOR(IO1I1OO00O1lIOOIll0lIO0l10lIlIIIII-1 DOWNTO 0);VARIABLE IO0Oll001000I1I0IIOO101lI10lIIIIII:STD_LOGIC_VECTOR(((4*II11OlI0I00OIO1llOI00O0lI0OlIIIIII)+7)-1 DOWNTO 0);VARIABLE
 IOI0IlOIlO11lO1OO1ll111101lO1IIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+2)-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE IIIlO001lO010I00O0OOllOO00l01IIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+2)-1 DOWNTO 0);VARIABLE IOlII0O0Oll1OO0O1O0O0O111O00lIIIII:
STD_LOGIC_VECTOR(IO0O010II00IOl10I10O1l0I10O1IOIIII DOWNTO 0);VARIABLE IOO1ll00l01O0lI100l10I1OOl0IIOIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+3)-1 DOWNTO 0);VARIABLE IO01Ol1OI1IO0OOIOIl01l001OI1OIIIII:STD_LOGIC_VECTOR(((2*IO0O010II00IOl10I10O1l0I10O1IOIIII)+5)-1
 DOWNTO 0);VARIABLE IOI111OlI111O1lI0lO1I00O0II10IIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+2)-1 DOWNTO 0);VARIABLE IIOI01II0OIl10O10OO010OIOllO0IIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+1)-1 DOWNTO 0);CONSTANT IOO0l1O1IlO1000Ol10IlOIO00111IIIII:
INTEGER:=(II1I1IOl0I0I1I0lIl00ll11I111OIIIII+IO0O010II00IOl10I10O1l0I10O1IOIIII+3);CONSTANT IOO0O01Il01I00O00IO0O0O1ll0O1IIIII:INTEGER:=(4*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3;VARIABLE IOOIl01IO0lllOIIlIO10l11I000lIIIII:STD_LOGIC_VECTOR(IOO0l1O1IlO1000Ol10IlOIO00111IIIII-1 DOWNTO 0):=(OTHERS
=>'0');VARIABLE III00lO01IIlOIllO00O0lIll1O1IIIIII:STD_LOGIC_VECTOR(IOO0l1O1IlO1000Ol10IlOIO00111IIIII-1 DOWNTO 0);CONSTANT IOlOI110lOlOI0OI11O000OOIl1IOIIIII:INTEGER:=IOO0l1O1IlO1000Ol10IlOIO00111IIIII-1-3-(IO0O010II00IOl10I10O1l0I10O1IOIIII-1);CONSTANT IO101lI0lO1OI00OIOO1lOI1l1lIIOIIII
:INTEGER:=IOO0l1O1IlO1000Ol10IlOIO00111IIIII-((4*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3);VARIABLE III11I1OOl0l0IIOIIIOOOIOl0010IIIII:STD_LOGIC_VECTOR((4*IO0O010II00IOl10I10O1l0I10O1IOIIII)-(IO0O010II00IOl10I10O1l0I10O1IOIIII-1)-1 DOWNTO 0);SUBTYPE IOlI00lO001l0IlOIOIlO11IOl011IIIII IS INTEGER RANGE III11I1OOl0l0IIOIIIOOOIOl0010IIIII'high DOWNTO
 III11I1OOl0l0IIOIIIOOOIOl0010IIIII'high+1-(IO0O010II00IOl10I10O1l0I10O1IOIIII+1);SUBTYPE IO1O0l0lO001lll1111lO1lOl100OIIIII IS INTEGER RANGE IOlI00lO001l0IlOIOIlO11IOl011IIIII'low-1 DOWNTO IOlI00lO001l0IlOIOIlO11IOl011IIIII'low-(IO0O010II00IOl10I10O1l0I10O1IOIIII);VARIABLE IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII:STD_LOGIC_VECTOR((IO0O010II00IOl10I10O1l0I10O1IOIIII+1)-1 DOWNTO
 0);VARIABLE IOIOlOOOOl01l0I1l0OI1Il1l1OO1IIIII:STD_LOGIC_VECTOR(IO0O010II00IOl10I10O1l0I10O1IOIIII-1 DOWNTO 0);VARIABLE IIlIIlIl01lOl1O00Ol00OOOIO1I0IIIII:STD_LOGIC_VECTOR(((2*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3)-1 DOWNTO 0):=(OTHERS=>'0');
VARIABLE II0I110I0IllOO1l11O1I0llOlOI1IIIII:STD_LOGIC_VECTOR(((2*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3)-1 DOWNTO 0);VARIABLE IOI1000Ol10O11I01I0O1lIII0OlIIIIII:STD_LOGIC_VECTOR(((3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+2)-1 DOWNTO 0);VARIABLE II1lOlIlO10lOOI0llO0lO1O0lO00IIIII:
STD_LOGIC_VECTOR(((3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3)-1 DOWNTO 0);VARIABLE IO0O100O1O0IlIl1OII1I0lOI0IO1IIIII:STD_LOGIC_VECTOR(((2*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3)-1 DOWNTO 0);VARIABLE II0I1O11I0IIlOlO111O1O0l010OIOIIII:STD_LOGIC_VECTOR(((3*IO0O010II00IOl10I10O1l0I10O1IOIIII
)+1)-1 DOWNTO 0);VARIABLE IOIOl1IO110100l0OIl0IIlIOO0IIOIIII:STD_LOGIC_VECTOR(((3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+2)-1 DOWNTO 0);VARIABLE III0ll0lIll1lIO11lOlIl0IO000IIIIII:STD_LOGIC_VECTOR(((5*IO0O010II00IOl10I10O1l0I10O1IOIIII)+2)-
1 DOWNTO 0);VARIABLE II10OIl0OO0IOIO111ll0Ill01l0OIIIII:STD_LOGIC_VECTOR(((5*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3)-1 DOWNTO 0);VARIABLE IIOlIIIIIlIIl0III10OO1OlI00lIOIIII:STD_LOGIC_VECTOR((II1I1IOl0I0I1I0lIl00ll11I111OIIIII-1)-1 DOWNTO 0);BEGIN IOI111lOI111OOlI0III1I0lO1I0IIIIII:=IOOl1IIO0I01ll0O00O01O1I000IOIIIII(IIOl00111100II1IOl0O1OO1I0lIOOIIII
+IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-1);II101I1OIIl111101l00ll0Ol1l01IIIII:=IOOl1IIO0I01ll0O00O01O1I000IOIIIII(IIOl00111100II1IOl0O1OO1I0lIOOIIII+IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-2 DOWNTO IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-1);IO1ll0OlO000O0lIO01I1llIOlOI1IIIII:=IOOl1IIO0I01ll0O00O01O1I000IOIIIII(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-2 DOWNTO 0);IOl0l0l0I0I0l0I010011l0llIl1lIIIII:=FLT_PT_IS_INF(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOOl1IIO0I01ll0O00O01O1I000IOIIIII);IO1l0OlOOl00O1OIlI0O0lIIlIlOlIIIII:=FLT_PT_IS_NAN(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOOl1IIO0I01ll0O00O01O1I000IOIIIII);II001lI100O0O0I1l1IIOlIlO00IlIIIII:=
II1IOOO1II0l1lOl00I1O001I00O0IIIII(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOOl1IIO0I01ll0O00O01O1I000IOIIIII);IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:='0';II0O01100OIIIl10O1OIl0I00Ol10IIIII:='0';IF IO1l0OlOOl00O1OIlI0O0lIIlIlOlIIIII THEN IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=FLT_PT_GET_QUIET_NAN(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII);ELSIF IOl0l0l0I0I0l0I010011l0llIl1lIIIII
 THEN IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=FLT_PT_GET_ZERO(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOI111lOI111OOlI0III1I0lO1I0IIIIII);ELSIF II001lI100O0O0I1l1IIOlIlO00IlIIIII THEN IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=FLT_PT_GET_INF(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOI111lOI111OOlI0III1I0lO1I0IIIIII);II0O01100OIIIl10O1OIl0I00Ol10IIIII:='1';ELSIF IO1ll0OlO000O0lIO01I1llIOlOI1IIIII=
FLT_PT_ZERO(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII-2 DOWNTO 0)THEN IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=IOI111lOI111OOlI0III1I0lO1I0IIIIII&STD_LOGIC_VECTOR(UNSIGNED(NOT(II101I1OIIl111101l00ll0Ol1l01IIIII))-TO_UNSIGNED(1,II101I1OIIl111101l00ll0Ol1l01IIIII'length))&IO1ll0OlO000O0lIO01I1llIOlOI1IIIII;IF TO_INTEGER(
UNSIGNED(NOT(II101I1OIIl111101l00ll0Ol1l01IIIII)))<=1 THEN IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:='1';ELSE IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:='0';END IF;ELSE IOOlII11IOO011lOll1IOO10O010OIIIII:=IO1ll0OlO000O0lIO01I1llIOlOI1IIIII(IO1ll0OlO000O0lIO01I1llIOlOI1IIIII'high DOWNTO IO1ll0OlO000O0lIO01I1llIOlOI1IIIII'high+1-IO0O010II00IOl10I10O1l0I10O1IOIIII);
IOI1IlOO001111I101I1O01l01lI1IIIII:=IOOlII11IOO011lOll1IOO10O010OIIIII(IO0O010II00IOl10I10O1l0I10O1IOIIII-1 DOWNTO IO0O010II00IOl10I10O1l0I10O1IOIIII-II11OlI0I00OIO1llOI00O0lI0OlIIIIII);II1l0l1O010I00O1Ill1O10lIII0OIIIII:=FLT_PT_RECIP_CALC_ROM_ENTRY(TO_INTEGER(UNSIGNED(IOI1IlOO001111I101I1O01l01lI1IIIII)),II11OlI0I00OIO1llOI00O0lI0OlIIIIII,IO1I1OO00O1lIOOIll0lIO0l10lIlIIIII);IO0Oll001000I1I0IIOO101lI10lIIIIII:=
STD_LOGIC_VECTOR(UNSIGNED(II1l0l1O010I00O1Ill1O10lIII0OIIIII)*UNSIGNED('1'&IOI1IlOO001111I101I1O01l01lI1IIIII&NOT(IOOlII11IOO011lOll1IOO10O010OIIIII(IO0O010II00IOl10I10O1l0I10O1IOIIII-II11OlI0I00OIO1llOI00O0lI0OlIIIIII-1 DOWNTO 0))&FLT_PT_ONE(((2*II11OlI0I00OIO1llOI00O0lI0OlIIIIII)-IO0O010II00IOl10I10O1l0I10O1IOIIII+3)-1 DOWNTO 0)));IOlII0O0Oll1OO0O1O0O0O111O00lIIIII:=IO0Oll001000I1I0IIOO101lI10lIIIIII(
IO0Oll001000I1I0IIOO101lI10lIIIIII'high-1 DOWNTO IO0Oll001000I1I0IIOO101lI10lIIIIII'high-(IO0O010II00IOl10I10O1l0I10O1IOIIII+1));IOO1ll00l01O0lI100l10I1OOl0IIOIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IOlII0O0Oll1OO0O1O0O0O111O00lIIIII)*UNSIGNED('1'&IOOlII11IOO011lOll1IOO10O010OIIIII),IO0O010II00IOl10I10O1l0I10O1IOIIII+3));IO01Ol1OI1IO0OOIOIl01l001OI1OIIIII:=
STD_LOGIC_VECTOR(-SIGNED(IOO1ll00l01O0lI100l10I1OOl0IIOIIII)*SIGNED('0'&IOlII0O0Oll1OO0O1O0O0O111O00lIIIII));IOI111OlI111O1lI0lO1I00O0II10IIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(IO01Ol1OI1IO0OOIOIl01l001OI1OIIIII(IO01Ol1OI1IO0OOIOIl01l001OI1OIIIII'high-1 DOWNTO IO01Ol1OI1IO0OOIOIl01l001OI1OIIIII'high
-3)),IO0O010II00IOl10I10O1l0I10O1IOIIII+2)+SIGNED('0'&IOlII0O0Oll1OO0O1O0O0O111O00lIIIII));IIOI01II0OIl10O10OO010OIOllO0IIIII:=IOI111OlI111O1lI0lO1I00O0II10IIIII(IOI111OlI111O1lI0lO1I00O0II10IIIII'high-1 DOWNTO 0);IOOIl01IO0lllOIIlIO10l11I000lIIIII(IOOIl01IO0lllOIIlIO10l11I000lIIIII'high DOWNTO IOOIl01IO0lllOIIlIO10l11I000lIIIII'high-2):=
"111";IOOIl01IO0lllOIIlIO10l11I000lIIIII(IOOIl01IO0lllOIIlIO10l11I000lIIIII'high-IOO0O01Il01I00O00IO0O0O1ll0O1IIIII):='1';III00lO01IIlOIllO00O0lIll1O1IIIIII:=STD_LOGIC_VECTOR(SIGNED(IOOIl01IO0lllOIIlIO10l11I000lIIIII)+(SIGNED(
'0'&IIOI01II0OIl10O10OO010OIOllO0IIIII)*SIGNED('0'&'1'&IO1ll0OlO000O0lIO01I1llIOlOI1IIIII)));III11I1OOl0l0IIOIIIOOOIOl0010IIIII:=III00lO01IIlOIllO00O0lIll1O1IIIIII(IOlOI110lOlOI0OI11O000OOIl1IOIIIII DOWNTO IO101lI0lO1OI00OIOO1lOI1l1lIIOIIII);IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII:=III11I1OOl0l0IIOIIIOOOIOl0010IIIII(IOlI00lO001l0IlOIOIlO11IOl011IIIII);IOIOlOOOOl01l0I1l0OI1Il1l1OO1IIIII:=III11I1OOl0l0IIOIIIOOOIOl0010IIIII(IO1O0l0lO001lll1111lO1lOl100OIIIII);IIlIIlIl01lOl1O00Ol00OOOIO1I0IIIII(0):='1'
;II0I110I0IllOO1l11O1I0llOlOI1IIIII:=STD_LOGIC_VECTOR(SIGNED(IIlIIlIl01lOl1O00Ol00OOOIO1I0IIIII)+(SIGNED(IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII)*SIGNED(IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII&'0')));IOI1000Ol10O11I01I0O1lIII0OlIIIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(II0I110I0IllOO1l11O1I0llOlOI1IIIII(II0I110I0IllOO1l11O1I0llOlOI1IIIII'high-1
 DOWNTO 0)&FLT_PT_ZERO((IO0O010II00IOl10I10O1l0I10O1IOIIII-1)-1 DOWNTO 0))+(SIGNED(IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII&'0')*SIGNED('0'&IOIOlOOOOl01l0I1l0OI1Il1l1OO1IIIII)),(3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+2));II1lOlIlO10lOOI0llO0lO1O0lO00IIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(IOI1000Ol10O11I01I0O1lIII0OlIIIIII)-(SIGNED
(II0I110I0IllOO1l11O1I0llOlOI1IIIII(II0I110I0IllOO1l11O1I0llOlOI1IIIII'high-1 DOWNTO II0I110I0IllOO1l11O1I0llOlOI1IIIII'high-(IO0O010II00IOl10I10O1l0I10O1IOIIII+1)))*SIGNED(IOIIOO0OlOOll0II1IOOI0IO0Il11IIIII)),(3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3));IO0O100O1O0IlIl1OII1I0lOI0IO1IIIII:=II1lOlIlO10lOOI0llO0lO1O0lO00IIIII(II1lOlIlO10lOOI0llO0lO1O0lO00IIIII'high DOWNTO II1lOlIlO10lOOI0llO0lO1O0lO00IIIII'high+1-((2*IO0O010II00IOl10I10O1l0I10O1IOIIII)+3));II0I1O11I0IIlOlO111O1O0l010OIOIIII:=III11I1OOl0l0IIOIIIOOOIOl0010IIIII(((3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+1
)-1 DOWNTO 0);IOIOl1IO110100l0OIl0IIlIOO0IIOIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(IO0O100O1O0IlIl1OII1I0lOI0IO1IIIII)-SIGNED(II0I1O11I0IIlOlO111O1O0l010OIOIIII),(3*IO0O010II00IOl10I10O1l0I10O1IOIIII)+2));III0ll0lIll1lIO11lOlIl0IO000IIIIII:='0'&IIOI01II0OIl10O10OO010OIOllO0IIIII&FLT_PT_ZERO((II1I1IOl0I0I1I0lIl00ll11I111OIIIII
-IO0O010II00IOl10I10O1l0I10O1IOIIII-1)-1 DOWNTO 0)&'1'&FLT_PT_ZERO(((4*IO0O010II00IOl10I10O1l0I10O1IOIIII)-II1I1IOl0I0I1I0lIl00ll11I111OIIIII+2+IO0O010II00IOl10I10O1l0I10O1IOIIII-2)-1 DOWNTO 0);II10OIl0OO0IOIO111ll0Ill01l0OIIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(III0ll0lIll1lIO11lOlIl0IO000IIIIII)+(
SIGNED('0'&IIOI01II0OIl10O10OO010OIOllO0IIIII)*SIGNED(IOIOl1IO110100l0OIl0IIlIOO0IIOIIII)),II10OIl0OO0IOIO111ll0Ill01l0OIIIII'length));IIOlIIIIIlIIl0III10OO1OlI00lIOIIII:=II10OIl0OO0IOIO111ll0Ill01l0OIIIII(II10OIl0OO0IOIO111ll0Ill01l0OIIIII'high-3 DOWNTO((5*IO0O010II00IOl10I10O1l0I10O1IOIIII)+1-II1I1IOl0I0I1I0lIl00ll11I111OIIIII));IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=IOI111lOI111OOlI0III1I0lO1I0IIIIII&STD_LOGIC_VECTOR(UNSIGNED(NOT(II101I1OIIl111101l00ll0Ol1l01IIIII
))-TO_UNSIGNED(2,II101I1OIIl111101l00ll0Ol1l01IIIII'length))&IIOlIIIIIlIIl0III10OO1OlI00lIOIIII;IF TO_INTEGER(UNSIGNED(NOT(II101I1OIIl111101l00ll0Ol1l01IIIII)))<=2 THEN IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:='1';ELSE IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII:='0';END IF;END
 IF;IF IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII='1'THEN IOO00I1Ill00Oll1OOOO01IlIlOlIIIIII:=FLT_PT_GET_ZERO(IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII+IIOl00111100II1IOl0O1OO1I0lIOOIIII,IOIII0l1O1IIOII0OI00lIOOI0IlOIIIII,IOI111lOI111OOlI0III1I0lO1I0IIIIII);END IF;III1lI0IOlOO11l0lO0IIl00OlOl0IIIII:=II0O01100OIIIl10O1OIl0I00Ol10IIIII;IIO1lIlIlIIll0011II00OlO00llOIIIII:=IOl0I1IOO010I0II10OOIl1ll1Ol1IIIII;END;
PROCEDURE IOll11O00IlllIl0l1I1I00l0IIOIIIIII(IIO1O11O1010OI0l1lI1IO0O1OlIIIIIII:IN INTEGER;IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII:IN INTEGER;IOI100O1O001OlIl001l1011IOll1IIIII:IN STD_LOGIC_VECTOR;IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:OUT STD_LOGIC_VECTOR;IOO0lIO01Ill01OO1Il00OO00I1l1IIIII:OUT STD_LOGIC
;IO11I0OIOIllIII10I01I1lO01IOIIIIII:OUT STD_LOGIC)IS CONSTANT IOIOll10I0lOl0I0IOOIl0IlI101IIIIII:INTEGER:=IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII;CONSTANT IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII:INTEGER:=IIO1O11O1010OI0l1lI1IO0O1OlIIIIIII-IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII;VARIABLE II0lO111OllO1OIl0IOlIIO011lllIIIII:STD_LOGIC_VECTOR(IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII-1 DOWNTO 0);
VARIABLE IOIIllIIII01O1l0OI1llO10Il1OIIIIII:STD_LOGIC_VECTOR(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO 0);VARIABLE IIO1llO1I11I00l1IIl1III0I0OOIOIIII:STD_LOGIC;VARIABLE IO1lllO01Il1110I10OIO0I01lIlOIIIII:BOOLEAN;VARIABLE II11llI1IOI1l1OI0I11ll1l1Ol0IOIIII:BOOLEAN;VARIABLE IOlIOIlOllOlO00IOO1I1IllIOll0IIIII:
BOOLEAN;VARIABLE IO11l0IlIIIlO10l0IlOI0OI1IOOlIIIII:STD_LOGIC_VECTOR(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII-1 DOWNTO 0);VARIABLE IIOOO001O1011l1OOO0I001lI0ll0IIIII:STD_LOGIC;VARIABLE IIIIOOI1OIl1IlOOI1OOOlIl0lOlIIIIII:STD_LOGIC;
CONSTANT II1I1l1lIIlO1lOOl10O0Oll100I0IIIII:INTEGER:=FLT_PT_RECIP_W(IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII);CONSTANT IOl0010llO1Ol00O0OOlII1I1IlI0IIIII:INTEGER:=FLT_PT_RECIP_K(IIO1O11O1010OI0l1lI1IO0O1OlIIIIIII,IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII,FLT_PT_RECIP_SQRT_OP_CODE);CONSTANT IO0O1II1OI11100IO0III1l1OI0IIIIIII:
INTEGER:=FLT_PT_RECIP_M(IIO1O11O1010OI0l1lI1IO0O1OlIIIIIII,IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII);CONSTANT IO0Ol000l0lOll0O0OOO0lOII00lIIIIII:INTEGER:=(2*IO0O1II1OI11100IO0III1l1OI0IIIIIII)+3;CONSTANT II1IIIlIl111lO10II01O1l0IOlIIIIIII:INTEGER:=(4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII);VARIABLE IOI0IIl1lIOI11l111I0I0lIIlOOlIIIII:
STD_LOGIC_VECTOR(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-1 DOWNTO 0);VARIABLE II01OOI10II1IIl1I11lI1II10IIOIIIII:STD_LOGIC_VECTOR(IO0O1II1OI11100IO0III1l1OI0IIIIIII-1 DOWNTO 0);VARIABLE IOlOlO1Illll100l0lO1OI11IIOllIIIII:STD_LOGIC_VECTOR(IO0Ol000l0lOll0O0OOO0lOII00lIIIIII-1
 DOWNTO 0);VARIABLE IIO0IIO0I000OIOIl1O00010Ill11IIIII:STD_LOGIC_VECTOR(((4*IO0O1II1OI11100IO0III1l1OI0IIIIIII)+7)-1 DOWNTO 0);VARIABLE II0IlOOIIlO0II0O1OOOIlOI1I10IIIIII:STD_LOGIC_VECTOR((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)-1 DOWNTO 0
):=(OTHERS=>'0');VARIABLE II1l1lO1IllI1OI1l0OlOOIl111OlIIIII:STD_LOGIC_VECTOR((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)-1 DOWNTO 0);VARIABLE IO0lIIllO0OIlIO0I1l0IIlII0l1IOIIII:STD_LOGIC_VECTOR(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII DOWNTO 0);VARIABLE IOlI1IlIO1O010Il1III1O0lO001IOIIII:
STD_LOGIC_VECTOR((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);VARIABLE IIlIl1100IO000lIO0l10IO1Ol01IOIIII:STD_LOGIC_VECTOR(((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)+5)-1 DOWNTO 0);VARIABLE IO0Il0OI0IOI0O1OIlO1I1IIO000lIIIII:STD_LOGIC_VECTOR((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)-1
 DOWNTO 0);VARIABLE IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII:STD_LOGIC_VECTOR((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE II1OO0I1Ill1I01lO1l0IllOlO11IIIIII:REAL;VARIABLE IOIOO1ll1O0Il0100001l1l1O1IIOOIIII:REAL;CONSTANT IO1lO0OOOI1111lOOl0lO00Il011IIIIII:REAL:=
REAL(1)/SQRT(REAL(2));VARIABLE IOII10010000l0II10OlOOllOl1IOIIIII:STD_LOGIC_VECTOR(II1IIIlIl111lO10II01O1l0IOlIIIIIII-1 DOWNTO 0);VARIABLE IOI1l0lII1II11Ill10III0111II1IIIII:STD_LOGIC_VECTOR(9 DOWNTO 0);VARIABLE
 IO1I01IOIlI0llO0OI0l10l00IlI0IIIII:REAL;VARIABLE IIll0O11I1IlIOOl1l100lOIOI1IIOIIII:SIGNED(17 DOWNTO 0);VARIABLE IO0Oll1llll1l100Il00OO110lO10IIIII:SIGNED(15 DOWNTO 0);VARIABLE III0IOl1OI0OO01O10OIlO0lO0OOIOIIII:SIGNED(35 DOWNTO 0);VARIABLE
 IO00l1llO0I0OOOI0II0I0O110111IIIII:SIGNED(35 DOWNTO 0);VARIABLE II1ll10l0OlO0OI0I1lOIIlOO1OOOIIIII:SIGNED(35 DOWNTO 0);VARIABLE IOIl11IO111IIl01O0lIlOlll01lIIIIII:SIGNED(24 DOWNTO 0);VARIABLE
 II11O1IllOlIO0I0l1IIIOIlO0l1OIIIII:SIGNED(40 DOWNTO 0);VARIABLE III1Ol01O00IO1ll0lO1OlIl1lO1lIIIII:SIGNED(40 DOWNTO 0);VARIABLE IIOlll0II1OlI00l10IlO0I1II101IIIII:SIGNED(40 DOWNTO 0);VARIABLE
 IIOl0Ollll00l0II0l0OO11O01ll1IIIII:SIGNED(24 DOWNTO 0);VARIABLE II0IIO1Ol0O1111I0OIOOOIIIOOO0IIIII:SIGNED(42 DOWNTO 0);VARIABLE IOO1IO1lIl1I0I00lO1lI0l1Ol1lOIIIII:SIGNED(34 DOWNTO 0);VARIABLE IOIOO11lIl00l11100lOI0llIIlO0IIIII:SIGNED
(69 DOWNTO 0);VARIABLE IIOl1OO0IOlIOll111O001lII1IlIIIIII:SIGNED(68 DOWNTO 0);VARIABLE IOlllIOI0IO1lIll001O0OlIOOIO0IIIII:SIGNED(84 DOWNTO 0);VARIABLE IOIII0IOl0O01O1IlII11O00lO101IIIII:SIGNED(84
 DOWNTO 0);VARIABLE II0ll0lI01OlIOl10lOO1I01OO0I1IIIII:SIGNED(84 DOWNTO 0);VARIABLE IOlIOOIIO01ll0lIlO1OIl001ll00IIIII:SIGNED(72 DOWNTO 0);VARIABLE IO1I1l0O00Oll0IO0llO0IOlI0O11IIIII:SIGNED(107 DOWNTO 0
);VARIABLE IOIOIOlOlOIIIII00OlI1OlIOOOlIOIIII:SIGNED(58 DOWNTO 0);VARIABLE IO1IOl10OlO0I00I00000O0l1O1OOIIIII:SIGNED(117 DOWNTO 0);VARIABLE IOllOII00lOI10lII1IIOI0OIl10lIIIII:SIGNED(117 DOWNTO 0);VARIABLE
 IO1IOlIl1lI1I1OllOI1Il1lI0Il1IIIII:SIGNED(117 DOWNTO 0);VARIABLE IOO01001IO0OO0lIIII1OII1I0lllIIIII:SIGNED(72 DOWNTO 0);VARIABLE III1O0l000IOIOIIOI1lIl11I01I0IIIII:SIGNED(88 DOWNTO 0);VARIABLE
 II0l0l1IO1lO111OI0I1lOO1lI1lIIIIII:SIGNED(88 DOWNTO 0);VARIABLE IIll0I0I1Il1l10Oll0lOI10OI0OlIIIII:SIGNED(88 DOWNTO 0);VARIABLE IOI1I011l1010IIll011lOO1I001OIIIII:SIGNED(58 DOWNTO 0);VARIABLE
 II10I1OIl1110OllIOllIIllI001IIIIII:SIGNED(117 DOWNTO 0);VARIABLE IOI0OO1l10I0l0l1l1OlI0O0IO01OIIIII:SIGNED(117 DOWNTO 0);VARIABLE IOIl0lI0I0I0Il11O0ll1lIlO00l1IIIII:SIGNED(117 DOWNTO 0);VARIABLE
 IOlO10l1OlIl1ll0IO1O1Il0I0I0OIIIII:SIGNED(58 DOWNTO 0);VARIABLE IIlllI1I1OOO1O0lI1I101010llO0IIIII:SIGNED(74 DOWNTO 0);VARIABLE III1OII01Ol1I01Ol1lO0O10110OIOIIII:SIGNED(74 DOWNTO 0);VARIABLE
 II0110IlI11OlIIO1IO1Il001100IOIIII:SIGNED(74 DOWNTO 0);VARIABLE IIOIlIO01Ol1O0l0I11l1OO1lOOO0IIIII:SIGNED(56 DOWNTO 0);CONSTANT IOOlOO01I10IllOlOIO0I0OllIOO0IIIII:UNSIGNED(55 DOWNTO 0
):=X"b504f333f9de65";CONSTANT IOl1l0I11OlI10Il10O1Ol10lI001IIIII:SIGNED(56 DOWNTO 0):=SIGNED(RESIZE(IOOlOO01I10IllOlOIO0I0OllIOO0IIIII,57));VARIABLE
 IOl0OOl01lIllOI0l1I00lO001lIIOIIII:SIGNED(113 DOWNTO 0);VARIABLE IIOlI1I0I0l0OlOI1OIIIIl1OlII1IIIII:SIGNED(113 DOWNTO 0);VARIABLE IIl0lIO0OO11l0O1OOlOO11OIOl0IOIIII:SIGNED(113 DOWNTO 0);
VARIABLE IOll1llllOOl1lIII11Il0OlO11llIIIII:SIGNED(56 DOWNTO 0);CONSTANT IIO1lOlIII0lIlOOI0ll011IO1I00IIIII:INTEGER:=(II1I1l1lIIlO1lOOl10O0Oll100I0IIIII+IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3);CONSTANT IO0lIIOO1Ol1l0OO10OIO010I1IIlIIIII:INTEGER:=(4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)+3;VARIABLE
 III11lO0lO1Ol0O10l001O11IIO01IIIII:STD_LOGIC_VECTOR(IIO1lOlIII0lIlOOI0ll011IO1I00IIIII-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE IIIOIl0O01O00OlIlIO0OIOII0O0lIIIII:STD_LOGIC_VECTOR(IIO1lOlIII0lIlOOI0ll011IO1I00IIIII-1 DOWNTO 0
);CONSTANT IO1lIOll10lIIOII1lI0Ill0O10IIOIIII:INTEGER:=IIO1lOlIII0lIlOOI0ll011IO1I00IIIII-1-3-(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-1);CONSTANT IOO0l1111I1l00OOOO0010l0OI001IIIII:INTEGER:=IIO1lOlIII0lIlOOI0ll011IO1I00IIIII-((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)+3);VARIABLE IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII:STD_LOGIC_VECTOR((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)-(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII
-1)-1 DOWNTO 0);SUBTYPE IO111010OOIOl0O1OIlIlI01010IOIIIII IS INTEGER RANGE IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII'high DOWNTO IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII'high+1-(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1);SUBTYPE II0II1l10O1OlI0Il000Ill10OOIOOIIII IS INTEGER RANGE IO111010OOIOl0O1OIlIlI01010IOIIIII'low-1
 DOWNTO IO111010OOIOl0O1OIlIlI01010IOIIIII'low-(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII);VARIABLE IO0O1l10lOlIO11Oll0OII00O0I0IIIIII:SIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IO010I000O1II100l01l0l1IlOOlOIIIII:UNSIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)-1 DOWNTO 0);VARIABLE IIOl1l0IO0O1lOI0I11l1I0llIOlOIIIII:SIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO
 0);VARIABLE IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII:SIGNED((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IIlllIlO1IIll0OIl1l0lllOI0OIIOIIII:SIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IOI10OlO11lI1011lI101Ol111I0IIIIII:SIGNED((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);
VARIABLE IIIl1I1O1llOllOO0OIO1l100I100IIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)-1 DOWNTO 0);VARIABLE IOO0l1IlO100O0II0IOI1l0O01I0OIIIII:SIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);VARIABLE IOl1IOlll1Il1Ol0l01I1001I1O0lIIIII:SIGNED((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+4)-1 DOWNTO 0
);VARIABLE IIOI0lll1IIO00lOl00I0OI1O11IIOIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);VARIABLE II01OIl1IOl11lO0OOO0lllIlI11IIIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+5)-1 DOWNTO 0);VARIABLE IOI11Il1OI0Illlll1l1OlII000OOIIIII:SIGNED((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+4)-1
 DOWNTO 0);VARIABLE II01IOI1OOO0I001Oll11I11OIlO0IIIII:SIGNED((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+5)-1 DOWNTO 0);VARIABLE IIII00IllI1lI1llI1011101OI0OOIIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+6)-1 DOWNTO 0);VARIABLE
 II1OlIO1IlO0000l00OIl1O111II1IIIII:SIGNED((2*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);VARIABLE IO1OO1IIIOl0llO0Ill11l1I00O10IIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IO1l001O0ll001lOl011I0O1lOI01IIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0);
VARIABLE IOllI1IO00I1II0OlO0OIl1ll01IlIIIII:SIGNED((3*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)-1 DOWNTO 0);VARIABLE IOOO0IlOO00ll1O0IOlO1IO0O11I0IIIII:STD_LOGIC_VECTOR((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IOl1I1010OOIlII1I1IOO00IOlIIIOIIII:STD_LOGIC_VECTOR
((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE II1OOl1OI0l1I1ll111110Ol1l00IOIIII:STD_LOGIC_VECTOR((8*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IIII0O0lO0ll110O1O1lIIOIOIII0IIIII:STD_LOGIC_VECTOR((7*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1
 DOWNTO 0);VARIABLE IO1I0001OI1l10O1lOO1l1l00l010IIIII:STD_LOGIC_VECTOR((8*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);VARIABLE IIOO10lOIllOOI101I0O0I1O10I1IOIIII:STD_LOGIC_VECTOR((8*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1)-1 DOWNTO 0);
VARIABLE IIl01OIlO0l1O0I010III11OO1IlIIIIII:STD_LOGIC_VECTOR((II1I1l1lIIlO1lOOl10O0Oll100I0IIIII-1)-1 DOWNTO 0);VARIABLE IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII:INTEGER;VARIABLE IOIl1OlI110lI10IO000lOIOIIO1lIIIII:STD_LOGIC_VECTOR(II0lO111OllO1OIl0IOlIIO011lllIIIII'range);
CONSTANT IO0010I1OOO1Ol1I1Il100001lIOlIIIII:INTEGER:=4*BOOLEAN'pos(FLT_PT_IS_DOUBLE_PRECISION(IIO1O11O1010OI0l1lI1IO0O1OlIIIIIII,IOl0OlI0OIlOIl11I0l0IlOOI01OOIIIII));BEGIN IIO1llO1I11I00l1IIl1III0I0OOIOIIII:=IOI100O1O001OlIl001l1011IOll1IIIII(IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII+IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-1);II0lO111OllO1OIl0IOlIIO011lllIIIII:=IOI100O1O001OlIl001l1011IOll1IIIII(IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII+IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO IOIOll10I0lOl0I0IOOIl0IlI101IIIIII
-1);IOIIllIIII01O1l0OI1llO10Il1OIIIIII:=IOI100O1O001OlIl001l1011IOll1IIIII(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO 0);IO1lllO01Il1110I10OIO0I01lIlOIIIII:=FLT_PT_IS_INF(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII,IOI100O1O001OlIl001l1011IOll1IIIII);II11llI1IOI1l1OI0I11ll1l1Ol0IOIIII:=FLT_PT_IS_NAN(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII,IOI100O1O001OlIl001l1011IOll1IIIII);IOlIOIlOllOlO00IOO1I1IllIOll0IIIII:=II1IOOO1II0l1lOl00I1O001I00O0IIIII(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII
,IOI100O1O001OlIl001l1011IOll1IIIII);IIOOO001O1011l1OOO0I001lI0ll0IIIII:='0';IIIIOOI1OIl1IlOOI1OOOlIl0lOlIIIIII:='0';IF II1I1l1lIIlO1lOOl10O0Oll100I0IIIII=24 THEN IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII:=127+(127/2);ELSE IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII:=1023+(1023/2);END IF;IF II11llI1IOI1l1OI0I11ll1l1Ol0IOIIII
 THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:=FLT_PT_GET_QUIET_NAN(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII);ELSIF IIO1llO1I11I00l1IIl1III0I0OOIOIIII='1'AND NOT(IOlIOIlOllOlO00IOO1I1IllIOll0IIIII)THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:=FLT_PT_GET_QUIET_NAN(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII);IIOOO001O1011l1OOO0I001lI0ll0IIIII:='1';ELSIF
 IO1lllO01Il1110I10OIO0I01lIlOIIIII THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:=FLT_PT_GET_ZERO(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII,IIO1llO1I11I00l1IIl1III0I0OOIOIIII);ELSIF IOlIOIlOllOlO00IOO1I1IllIOll0IIIII THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:=FLT_PT_GET_INF(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII+IOl0OO0lOI1O0l0I1lIlI00lO0llOIIIII,IOIOll10I0lOl0I0IOOIl0IlI101IIIIII,IIO1llO1I11I00l1IIl1III0I0OOIOIIII);IIIIOOI1OIl1IlOOI1OOOlIl0lOlIIIIII:='1';ELSIF IOIIllIIII01O1l0OI1llO10Il1OIIIIII=
FLT_PT_ZERO(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO 0)THEN IOIl1OlI110lI10IO000lOIOIIO1lIIIII:=STD_LOGIC_VECTOR(UNSIGNED(II0lO111OllO1OIl0IOlIIO011lllIIIII)SRL 1);IF II0lO111OllO1OIl0IOlIIO011lllIIIII(0)='1'THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:='0'&STD_LOGIC_VECTOR(
TO_UNSIGNED(IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII,II0lO111OllO1OIl0IOlIIO011lllIIIII'length)-UNSIGNED(IOIl1OlI110lI10IO000lOIOIIO1lIIIII))&IOIIllIIII01O1l0OI1llO10Il1OIIIIII;ELSE IF II1I1l1lIIlO1lOOl10O0Oll100I0IIIII=24 THEN IOIIllIIII01O1l0OI1llO10Il1OIIIIII:=FLT_PT_SQRT2_SGL(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO 0);ELSE
 IOIIllIIII01O1l0OI1llO10Il1OIIIIII:=FLT_PT_SQRT2_DBL(IOIOll10I0lOl0I0IOOIl0IlI101IIIIII-2 DOWNTO 0);END IF;IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:='0'&STD_LOGIC_VECTOR(TO_UNSIGNED(IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII,II0lO111OllO1OIl0IOlIIO011lllIIIII'length)-UNSIGNED(
IOIl1OlI110lI10IO000lOIOIIO1lIIIII))&IOIIllIIII01O1l0OI1llO10Il1OIIIIII;END IF;ELSE IOI0IIl1lIOI11l111I0I0lIIlOOlIIIII:=IOIIllIIII01O1l0OI1llO10Il1OIIIIII(IOIIllIIII01O1l0OI1llO10Il1OIIIIII'high DOWNTO IOIIllIIII01O1l0OI1llO10Il1OIIIIII'high+1-IOl0010llO1Ol00O0OOlII1I1IlI0IIIII);II01OOI10II1IIl1I11lI1II10IIOIIIII:=IOI0IIl1lIOI11l111I0I0lIIlOOlIIIII(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-1 DOWNTO IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-IO0O1II1OI11100IO0III1l1OI0IIIIIII);IOlOlO1Illll100l0lO1OI11IIOllIIIII:=
FLT_PT_RECIP_CALC_ROM_ENTRY(TO_INTEGER(UNSIGNED(II01OOI10II1IIl1I11lI1II10IIOIIIII)),IO0O1II1OI11100IO0III1l1OI0IIIIIII,IO0Ol000l0lOll0O0OOO0lOII00lIIIIII);IIO0IIO0I000OIOIl1O00010Ill11IIIII:=STD_LOGIC_VECTOR(UNSIGNED(IOlOlO1Illll100l0lO1OI11IIOllIIIII)*
UNSIGNED('1'&II01OOI10II1IIl1I11lI1II10IIOIIIII&NOT(IOI0IIl1lIOI11l111I0I0lIIlOOlIIIII(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-IO0O1II1OI11100IO0III1l1OI0IIIIIII-1 DOWNTO 0))&FLT_PT_ONE(((2*IO0O1II1OI11100IO0III1l1OI0IIIIIII)-IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3)-1 DOWNTO 0)));IO0lIIllO0OIlIO0I1l0IIlII0l1IOIIII:=IIO0IIO0I000OIOIl1O00010Ill11IIIII(IIO0IIO0I000OIOIl1O00010Ill11IIIII'high-1 DOWNTO
 IIO0IIO0I000OIOIl1O00010Ill11IIIII'high-(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1));IOlI1IlIO1O010Il1III1O0lO001IOIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IO0lIIllO0OIlIO0I1l0IIlII0l1IOIIII)*UNSIGNED('1'&IOI0IIl1lIOI11l111I0I0lIIlOOlIIIII),IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+3));IIlIl1100IO000lIO0l10IO1Ol01IOIIII:=STD_LOGIC_VECTOR(-SIGNED(
IOlI1IlIO1O010Il1III1O0lO001IOIIII)*SIGNED('0'&IO0lIIllO0OIlIO0I1l0IIlII0l1IOIIII));IO0Il0OI0IOI0O1OIlO1I1IIO000lIIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(IIlIl1100IO000lIO0l10IO1Ol01IOIIII(IIlIl1100IO000lIO0l10IO1Ol01IOIIII'high-1 DOWNTO IIlIl1100IO000lIO0l10IO1Ol01IOIIII'high-3)),IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+2)+SIGNED('0'&
IO0lIIllO0OIlIO0I1l0IIlII0l1IOIIII));IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII:=IO0Il0OI0IOI0O1OIlO1I1IIO000lIIIII(IO0Il0OI0IOI0O1OIlO1I1IIO000lIIIII'high-1 DOWNTO 0);III11lO0lO1Ol0O10l001O11IIO01IIIII(III11lO0lO1Ol0O10l001O11IIO01IIIII'high DOWNTO III11lO0lO1Ol0O10l001O11IIO01IIIII'high-2):="111";III11lO0lO1Ol0O10l001O11IIO01IIIII(
III11lO0lO1Ol0O10l001O11IIO01IIIII'high-IO0lIIOO1Ol1l0OO10OIO010I1IIlIIIII):='1';IIIOIl0O01O00OlIlIO0OIOII0O0lIIIII:=STD_LOGIC_VECTOR(SIGNED(III11lO0lO1Ol0O10l001O11IIO01IIIII)+(SIGNED('0'&IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII)*SIGNED('0'&'1'&
IOIIllIIII01O1l0OI1llO10Il1OIIIIII)));IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII:=IIIOIl0O01O00OlIlIO0OIOII0O0lIIIII(IO1lIOll10lIIOII1lI0Ill0O10IIOIIII DOWNTO IOO0l1111I1l00OOOO0010l0OI001IIIII);IF II1I1l1lIIlO1lOOl10O0Oll100I0IIIII=24 THEN II1OO0I1Ill1I01lO1l0IllOlO11IIIIII:=REAL(TO_INTEGER(UNSIGNED(IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII)))/REAL(2)**(IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1);IOIOO1ll1O0Il0100001l1l1O1IIOOIIII:=SQRT
(II1OO0I1Ill1I01lO1l0IllOlO11IIIIII);IF II0lO111OllO1OIl0IOlIIO011lllIIIII(0)='0'THEN IOII10010000l0II10OlOOllOl1IOIIIII:=STD_LOGIC_VECTOR(RESIZE(TO_UNSIGNED(INTEGER(ROUND(IOIOO1ll1O0Il0100001l1l1O1IIOOIIII*IO1lO0OOOI1111lOOl0lO00Il011IIIIII*REAL(2)**(4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII))),II1IIIlIl111lO10II01O1l0IOlIIIIIII),
II1IIIlIl111lO10II01O1l0IOlIIIIIII));ELSE IOII10010000l0II10OlOOllOl1IOIIIII:=STD_LOGIC_VECTOR(RESIZE(TO_UNSIGNED(INTEGER(ROUND(IOIOO1ll1O0Il0100001l1l1O1IIOOIIII*REAL(2)**(4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII))),II1IIIlIl111lO10II01O1l0IOlIIIIIII),II1IIIlIl111lO10II01O1l0IOlIIIIIII));END IF;ELSE IOI1l0lII1II11Ill10III0111II1IIIII
:=IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII(IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII'high DOWNTO IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII'high-9);II1OO0I1Ill1I01lO1l0IllOlO11IIIIII:=(REAL(TO_INTEGER(UNSIGNED(IOI1l0lII1II11Ill10III0111II1IIIII)))+REAL(1))/REAL(2)**10;IOIOO1ll1O0Il0100001l1l1O1IIOOIIII:=CEIL(SQRT(II1OO0I1Ill1I01lO1l0IllOlO11IIIIII)*REAL(2)**34
)/REAL(2)**34;IO1I01IOIlI0llO0OI0l10l00IlI0IIIII:=REAL(1)/IOIOO1ll1O0Il0100001l1l1O1IIOOIIII;IIll0O11I1IlIOOl1l100lOIOI1IIOIIII:=TO_SIGNED(INTEGER(FLOOR(IO1I01IOIlI0llO0OI0l10l00IlI0IIIII*REAL(2)**16)),18);IO0Oll1llll1l100Il00OO110lO10IIIII:=SIGNED(RESIZE(UNSIGNED(IOI0l1OOO0lllllI1l1OIOO0I1Il1IIIII),16));
III0IOl1OI0OO01O10OIlO0lO0OOIOIIII:=IIll0O11I1IlIOOl1l100lOIOI1IIOIIII*IIll0O11I1IlIOOl1l100lOIOI1IIOIIII;IO00l1llO0I0OOOI0II0I0O110111IIIII:=(9=>'1',OTHERS=>'0');II1ll10l0OlO0OI0I1lOIIlOO1OOOIIIII:=III0IOl1OI0OO01O10OIlO0lO0OOIOIIII+IO00l1llO0I0OOOI0II0I0O110111IIIII;IOIl11IO111IIl01O0lIlOlll01lIIIIII:=II1ll10l0OlO0OI0I1lOIIlOO1OOOIIIII(34 DOWNTO
 10);II11O1IllOlIO0I0l1IIIOIlO0l1OIIIII:=IO0Oll1llll1l100Il00OO110lO10IIIII*IOIl11IO111IIl01O0lIlOlll01lIIIIII;III1Ol01O00IO1ll0lO1OlIl1lO1lIIIII:=(38=>'1',37=>'1',14=>'1',OTHERS=>'0');IIOlll0II1OlI00l10IlO0I1II101IIIII:=III1Ol01O00IO1ll0lO1OlIl1lO1lIIIII-II11O1IllOlIO0I0l1IIIOIlO0l1OIIIII;
IIOl0Ollll00l0II0l0OO11O01ll1IIIII:=IIOlll0II1OlI00l10IlO0I1II101IIIII(39 DOWNTO 15);II0IIO1Ol0O1111I0OIOOOIIIOOO0IIIII:=IIll0O11I1IlIOOl1l100lOIOI1IIOIIII*IIOl0Ollll00l0II0l0OO11O01ll1IIIII;IOO1IO1lIl1I0I00lO1lI0l1Ol1lOIIIII:=II0IIO1Ol0O1111I0OIOOOIIIOOO0IIIII(40 DOWNTO 6);IOIOO11lIl00l11100lOI0llIIlO0IIIII:=IOO1IO1lIl1I0I00lO1lI0l1Ol1lOIIIII*IOO1IO1lIl1I0I00lO1lI0l1Ol1lOIIIII;IIOl1OO0IOlIOll111O001lII1IlIIIIII:=IOIOO11lIl00l11100lOI0llIIlO0IIIII
(68 DOWNTO 0);IOlllIOI0IO1lIll001O0OlIOOIO0IIIII:=IO0Oll1llll1l100Il00OO110lO10IIIII*IIOl1OO0IOlIOll111O001lII1IlIIIIII;IOIII0IOl0O01O1IlII11O00lO101IIIII:=(82=>'1',81=>'1',10=>'1',OTHERS=>'0');II0ll0lI01OlIOl10lOO1I01OO0I1IIIII:=IOIII0IOl0O01O1IlII11O00lO101IIIII-
IOlllIOI0IO1lIll001O0OlIOOIO0IIIII;IOlIOOIIO01ll0lIlO1OIl001ll00IIIII:=II0ll0lI01OlIOl10lOO1I01OO0I1IIIII(83 DOWNTO 11);IO1I1l0O00Oll0IO0llO0IOlI0O11IIIII:=IOO1IO1lIl1I0I00lO1lI0l1Ol1lOIIIII*IOlIOOIIO01ll0lIlO1OIl001ll00IIIII;IOIOIOlOlOIIIII00OlI1OlIOOOlIOIIII:=IO1I1l0O00Oll0IO0llO0IOlI0O11IIIII(105 DOWNTO 47);IO1IOl10OlO0I00I00000O0l1O1OOIIIII:=IOIOIOlOlOIIIII00OlI1OlIOOOlIOIIII*IOIOIOlOlOIIIII00OlI1OlIOOOlIOIIII;
IOllOII00lOI10lII1IIOI0OIl10lIIIII:=(43=>'1',OTHERS=>'0');IO1IOlIl1lI1I1OllOI1Il1lI0Il1IIIII:=IO1IOl10OlO0I00I00000O0l1O1OOIIIII+IOllOII00lOI10lII1IIOI0OIl10lIIIII;IOO01001IO0OO0lIIII1OII1I0lllIIIII:=IO1IOlIl1lI1I1OllOI1Il1lI0Il1IIIII(116 DOWNTO 44);III1O0l000IOIOIIOI1lIl11I01I0IIIII:=
IO0Oll1llll1l100Il00OO110lO10IIIII*IOO01001IO0OO0lIIII1OII1I0lllIIIII;II0l0l1IO1lO111OI0I1lOO1lI1lIIIIII:=(86=>'1',85=>'1',28=>'1',OTHERS=>'0');IIll0I0I1Il1l10Oll0lOI10OI0OlIIIII:=II0l0l1IO1lO111OI0I1lOO1lI1lIIIIII-III1O0l000IOIOIIOI1lIl11I01I0IIIII;IOI1I011l1010IIll011lOO1I001OIIIII:=IIll0I0I1Il1l10Oll0lOI10OI0OlIIIII(
87 DOWNTO 29);II10I1OIl1110OllIOllIIllI001IIIIII:=IOIOIOlOlOIIIII00OlI1OlIOOOlIOIIII*IOI1I011l1010IIll011lOO1I001OIIIII;IOI0OO1l10I0l0l1l1OlI0O0IO01OIIIII:=(56=>'1',OTHERS=>'0');IOIl0lI0I0I0Il11O0ll1lIlO00l1IIIII:=II10I1OIl1110OllIOllIIllI001IIIIII+IOI0OO1l10I0l0l1l1OlI0O0IO01OIIIII;IOlO10l1OlIl1ll0IO1O1Il0I0I0OIIIII:=
IOIl0lI0I0I0Il11O0ll1lIlO00l1IIIII(115 DOWNTO 57);IIlllI1I1OOO1O0lI1I101010llO0IIIII:=IOlO10l1OlIl1ll0IO1O1Il0I0I0OIIIII*IO0Oll1llll1l100Il00OO110lO10IIIII;III1OII01Ol1I01Ol1lO0O10110OIOIIII:=(15=>'1',OTHERS=>'0');II0110IlI11OlIIO1IO1Il001100IOIIII:=IIlllI1I1OOO1O0lI1I101010llO0IIIII
+III1OII01Ol1I01Ol1lO0O10110OIOIIII;IIOIlIO01Ol1O0l0I11l1OO1lOOO0IIIII:=II0110IlI11OlIIO1IO1Il001100IOIIII(72 DOWNTO 16);IF II0lO111OllO1OIl0IOlIIO011lllIIIII(0)='0'THEN IOl0OOl01lIllOI0l1I00lO001lIIOIIII:=IIOIlIO01Ol1O0l0I11l1OO1lOOO0IIIII*
IOl1l0I11OlI10Il10O1Ol10lI001IIIII;IIOlI1I0I0l0OlOI1OIIIIl1OlII1IIIII:=(55=>'1',OTHERS=>'0');IIl0lIO0OO11l0O1OOlOO11OIOl0IOIIII:=IOl0OOl01lIllOI0l1I00lO001lIIOIIII+IIOlI1I0I0l0OlOI1OIIIIl1OlII1IIIII;IOll1llllOOl1lIII11Il0OlO11llIIIII:=IIl0lIO0OO11l0O1OOlOO11OIOl0IOIIII
(112 DOWNTO 56);ELSE IOll1llllOOl1lIII11Il0OlO11llIIIII:=IIOIlIO01Ol1O0l0I11l1OO1lOOO0IIIII;END IF;IOII10010000l0II10OlOOllOl1IOIIIII:=STD_LOGIC_VECTOR(RESIZE(UNSIGNED(IOll1llllOOl1lIII11Il0OlO11llIIIII),II1IIIlIl111lO10II01O1l0IOlIIIIIII));END IF;IO0O1l10lOlIO11Oll0OII00O0I0IIIIII:=SIGNED(IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII(
IO111010OOIOl0O1OIlIlI01010IOIIIII));IO010I000O1II100l01l0l1IlOOlOIIIII:=UNSIGNED(IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII(II0II1l10O1OlI0Il000Ill10OOIOOIIII));IIOl1l0IO0O1lOI0I11l1I0llIOlOIIIII:=SIGNED(RESIZE(IO010I000O1II100l01l0l1IlOOlOIIIII,IIOl1l0IO0O1lOI0I11l1I0llIOlOIIIII'length));IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII:=RESIZE(IO0O1l10lOlIO11Oll0OII00O0I0IIIIII*IO0O1l10lOlIO11Oll0OII00O0I0IIIIII,IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII'length);IIlllIlO1IIll0OIl1l0lllOI0OIIOIIII:=IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII(IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII'high DOWNTO IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII
'high-IIlllIlO1IIll0OIl1l0lllOI0OIIOIIII'length+1);IOI10OlO11lI1011lI101Ol111I0IIIIII:=RESIZE(IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII,IOI10OlO11lI1011lI101Ol111I0IIIIII'length)+RESIZE(IO1l1l0O010OlO0I1ll1O1lI1I0I1IIIII&'0',IOI10OlO11lI1011lI101Ol111I0IIIIII'length);IIIl1I1O1llOllOO0OIO1l100I100IIIII:=IOI10OlO11lI1011lI101Ol111I0IIIIII&SIGNED(FLT_PT_ZERO((IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-1)-1
 DOWNTO 0));IOO0l1IlO100O0II0IOI1l0O01I0OIIIII:=RESIZE(IIOl1l0IO0O1lOI0I11l1I0llIOlOIIIII,IOO0l1IlO100O0II0IOI1l0O01I0OIIIII'length)+RESIZE(IIOl1l0IO0O1lOI0I11l1I0llIOlOIIIII&'0',IOO0l1IlO100O0II0IOI1l0O01I0OIIIII'length);IOl1IOlll1Il1Ol0l01I1001I1O0lIIIII:=IOO0l1IlO100O0II0IOI1l0O01I0OIIIII*IO0O1l10lOlIO11Oll0OII00O0I0IIIIII;IIOI0lll1IIO00lOl00I0OI1O11IIOIIII:=RESIZE(IOl1IOlll1Il1Ol0l01I1001I1O0lIIIII,IIOI0lll1IIO00lOl00I0OI1O11IIOIIII'length
)+RESIZE(IIIl1I1O1llOllOO0OIO1l100I100IIIII,IIOI0lll1IIO00lOl00I0OI1O11IIOIIII'length);II01OIl1IOl11lO0OOO0lllIlI11IIIIII:=IIOI0lll1IIO00lOl00I0OI1O11IIOIIII&"00";IOI11Il1OI0Illlll1l1OlII000OOIIIII:=RESIZE(IO0O1l10lOlIO11Oll0OII00O0I0IIIIII,IOI11Il1OI0Illlll1l1OlII000OOIIIII'length)+RESIZE(IO0O1l10lOlIO11Oll0OII00O0I0IIIIII&"00",IOI11Il1OI0Illlll1l1OlII000OOIIIII'length);
II01IOI1OOO0I001Oll11I11OIlO0IIIII:=IIlllIlO1IIll0OIl1l0lllOI0OIIOIIII*IOI11Il1OI0Illlll1l1OlII000OOIIIII;IIII00IllI1lI1llI1011101OI0OOIIIII:=RESIZE(II01OIl1IOl11lO0OOO0lllIlI11IIIIII,IIII00IllI1lI1llI1011101OI0OOIIIII'length)-RESIZE(II01IOI1OOO0I001Oll11I11OIlO0IIIII,IIII00IllI1lI1llI1011101OI0OOIIIII'length);
II1OlIO1IlO0000l00OIl1O111II1IIIII:=IIII00IllI1lI1llI1011101OI0OOIIIII(IIII00IllI1lI1llI1011101OI0OOIIIII'high DOWNTO IIII00IllI1lI1llI1011101OI0OOIIIII'high-II1OlIO1IlO0000l00OIl1O111II1IIIII'length+1);IO1OO1IIIOl0llO0Ill11l1I00O10IIIII:=SIGNED(IIOIOl1l11I0OO0l1OO1llIOIllO0IIIII);IO1l001O0ll001lOl011I0O1lOI01IIIII:=RESIZE
(II1OlIO1IlO0000l00OIl1O111II1IIIII,IO1l001O0ll001lOl011I0O1lOI01IIIII'length)-RESIZE(IO1OO1IIIOl0llO0Ill11l1I00O10IIIII,IO1l001O0ll001lOl011I0O1lOI01IIIII'length)+TO_SIGNED(1,IO1l001O0ll001lOl011I0O1lOI01IIIII'length);IOllI1IO00I1II0OlO0OIl1ll01IlIIIII:=IO1l001O0ll001lOl011I0O1lOI01IIIII(IO1l001O0ll001lOl011I0O1lOI01IIIII'high DOWNTO 1);IOOO0IlOO00ll1O0IOlO1IO0O11I0IIIII
:=FLT_PT_ZERO((II1I1l1lIIlO1lOOl10O0Oll100I0IIIII+1)-1 DOWNTO 0)&'1'&FLT_PT_ZERO((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII-II1I1l1lIIlO1lOOl10O0Oll100I0IIIII-1)-1 DOWNTO 0);IOl1I1010OOIlII1I1IOO00IOlIIIOIIII:=STD_LOGIC_VECTOR(SIGNED('0'&IOII10010000l0II10OlOOllOl1IOIIIII)+SIGNED(IOOO0IlOO00ll1O0IOlO1IO0O11I0IIIII))
;IIII0O0lO0ll110O1O1lIIOIOIII0IIIII:=STD_LOGIC_VECTOR(SIGNED('0'&IOII10010000l0II10OlOOllOl1IOIIIII)*SIGNED(IOllI1IO00I1II0OlO0OIl1ll01IlIIIII));IO1I0001OI1l10O1lOO1l1l00l010IIIII:=STD_LOGIC_VECTOR(RESIZE(SIGNED(IIII0O0lO0ll110O1O1lIIOIOIII0IIIII),8*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII+1));
II1OOl1OI0l1I1ll111110Ol1l00IOIIII:=IOl1I1010OOIlII1I1IOO00IOlIIIOIIII&FLT_PT_ZERO((4*IOl0010llO1Ol00O0OOlII1I1IlI0IIIII)-1 DOWNTO 0);IIOO10lOIllOOI101I0O0I1O10I1IOIIII:=STD_LOGIC_VECTOR(SIGNED(IO1I0001OI1l10O1lOO1l1l00l010IIIII)+SIGNED(
II1OOl1OI0l1I1ll111110Ol1l00IOIIII));IIl01OIlO0l1O0I010III11OO1IlIIIIII:=IIOO10lOIllOOI101I0O0I1O10I1IOIIII(IIOO10lOIllOOI101I0O0I1O10I1IOIIII'high-2 DOWNTO IIOO10lOIllOOI101I0O0I1O10I1IOIIII'high-II1I1l1lIIlO1lOOl10O0Oll100I0IIIII);IOIl1OlI110lI10IO000lOIOIIO1lIIIII:=STD_LOGIC_VECTOR(UNSIGNED(II0lO111OllO1OIl0IOlIIO011lllIIIII)SRL 1);IF II0lO111OllO1OIl0IOlIIO011lllIIIII
(0)='1'THEN IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:='0'&STD_LOGIC_VECTOR(TO_UNSIGNED(IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII-1,II0lO111OllO1OIl0IOlIIO011lllIIIII'length)-UNSIGNED(IOIl1OlI110lI10IO000lOIOIIO1lIIIII))&IIl01OIlO0l1O0I010III11OO1IlIIIIII;ELSE IO0l1OlI0l011l0lO1O11OlOO0lllIIIII:='0'&
STD_LOGIC_VECTOR(TO_UNSIGNED(IOO00OI01Ol1l0lIlOO1lI0OI11I0IIIII,II0lO111OllO1OIl0IOlIIO011lllIIIII'length)-UNSIGNED(IOIl1OlI110lI10IO000lOIOIIO1lIIIII))&IIl01OIlO0l1O0I010III11OO1IlIIIIII;END IF;END IF;IOO0lIO01Ill01OO1Il00OO00I1l1IIIII:=IIIIOOI1OIl1IlOOI1OOOlIl0lOlIIIIII;
IO11I0OIOIllIII10I01I1lO01IOIIIIII:=IIOOO001O1011l1OOO0I001lI0ll0IIIII;END;PROCEDURE II11l0O1IO1OOI000IIO11I1Oll1IIIIII(IOO011IOl1001I1O1lIOOIlO0l01IIIIII:IN STD_LOGIC_VECTOR(C_A_WIDTH-1 DOWNTO 0);IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII:IN STD_LOGIC_VECTOR(C_B_WIDTH-1
 DOWNTO 0);IOlOII1IIOlI01OI0IOOIllI0I1IOIIIII:IN STD_LOGIC_VECTOR(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0);IOOl0O0Il1Il00ll0l0l110I1OIllIIIII:OUT STD_LOGIC_VECTOR(C_RESULT_WIDTH-1 DOWNTO 0);
IIO0lO00IO0IO01O001OIOlll11OlIIIII:OUT STD_LOGIC;II000llI0IIOIlO0OO01I11I01000IIIII:OUT STD_LOGIC;II1IIlIllI0l0O110Il0OlIII1OOOIIIII:OUT STD_LOGIC;IIO0ll0III00OIOOI1I1OI1lIlO1OIIIII:OUT STD_LOGIC)IS VARIABLE IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII:
STD_LOGIC_VECTOR(C_RESULT_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE IO0010l0I011lIOIOOl1O1l101lllIIIII:STD_LOGIC;VARIABLE IOOOOOl1OOO010IO00O0IO0Il10O1IIIII:STD_LOGIC;
VARIABLE IOllIl0O0Ollll0IOlI011lI01Il1IIIII:STD_LOGIC;VARIABLE IO1IOI00OI0I10OO1l0I0l1l010llIIIII:STD_LOGIC;VARIABLE IO10I111l1OOlIO0IlI1I00llll0lIIIII:BOOLEAN;BEGIN IO0010l0I011lIOIOOl1O1l101lllIIIII:='0';
IOOOOOl1OOO010IO00O0IO0Il10O1IIIII:='0';IOllIl0O0Ollll0IOlI011lI01Il1IIIII:='0';IO1IOI00OI0I10OO1l0I0l1l010llIIIII:='0';IO10I111l1OOlIO0IlI1I00llll0lIIIII:=FALSE;CASE TO_INTEGER(UNSIGNED(IOlOII1IIOlI01OI0IOOIllI0I1IOIIIII(FLT_PT_OP_CODE_SLICE)))
IS WHEN FLT_PT_SQRT_OP_CODE=>IF(C_HAS_SQRT=FLT_PT_YES)THEN IF((C_RESULT_WIDTH=C_A_WIDTH)AND(C_RESULT_FRACTION_WIDTH=
C_A_FRACTION_WIDTH))THEN IOOll1I1OOlO0lOO0IIII1lO11IIlIIIII(C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);
IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;ELSIF(C_HAS_FLT_TO_FLT=FLT_PT_YES)THEN IO1I1OlOI1OII110llI1lI0IIl0O0IIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,C_RESULT_WIDTH,
C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;ELSIF(C_HAS_RECIP=FLT_PT_YES)THEN
 IF((C_RESULT_WIDTH=C_A_WIDTH)AND(C_RESULT_FRACTION_WIDTH=C_A_FRACTION_WIDTH))THEN IOOOOI1lIlOlI10IOOOI00O10O00IIIIII(C_RESULT_WIDTH,
C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IOllIl0O0Ollll0IOlI011lI01Il1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;ELSIF(C_HAS_RECIP_SQRT=FLT_PT_YES)
THEN IF((C_RESULT_WIDTH=C_A_WIDTH)AND(C_RESULT_FRACTION_WIDTH=C_A_FRACTION_WIDTH))THEN IOll11O00IlllIl0l1I1I00l0IIOIIIIII(C_RESULT_WIDTH,
C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IOllIl0O0Ollll0IOlI011lI01Il1IIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;END IF;WHEN FLT_PT_DIVIDE_OP_CODE
=>IF(C_HAS_DIVIDE=FLT_PT_YES)THEN II1lIII001001Il0l0OOl0I00I01IIIIII(C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,
IO1IOI00OI0I10OO1l0I0l1l010llIIIII,IOllIl0O0Ollll0IOlI011lI01Il1IIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;WHEN FLT_PT_MULTIPLY_OP_CODE=>IF(C_HAS_MULTIPLY=FLT_PT_YES)THEN
 IIOOO0OOIll110IlI1111I1001I01IIIII(C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE
;END IF;WHEN FLT_PT_ADD_OP_CODE=>IF C_HAS_ADD=FLT_PT_TRUE THEN IOO0llOIlIO0110l1lOO01I00l1OIIIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,FALSE,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,
IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;WHEN FLT_PT_SUBTRACT_OP_CODE=>IF C_HAS_SUBTRACT=FLT_PT_TRUE
 THEN IOO0llOIlIO0110l1lOO01I00l1OIIIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,TRUE,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END
 IF;WHEN FLT_PT_COMPARE_OP_CODE=>IF(C_HAS_COMPARE=FLT_PT_YES)THEN IO1lII1OIl0llIl0IIlIlOI10l0OlIIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,C_RESULT_WIDTH,IOlOII1IIOlI01OI0IOOIllI0I1IOIIIII(
FLT_PT_COMPARE_OPERATION_SLICE),IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;WHEN FLT_PT_FLT_TO_FIX_OP_CODE=>IF(
C_HAS_FLT_TO_FIX=FLT_PT_YES)THEN II1011l1lI11IlIlI0l0l00100lO0IIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII
,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;WHEN FLT_PT_FIX_TO_FLT_OP_CODE=>IF(C_HAS_FIX_TO_FLT=FLT_PT_YES
)THEN II111O1llOOlI0lOOIIIl0OIlIlllIIIII(C_A_WIDTH,C_A_FRACTION_WIDTH,C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH,IOO011IOl1001I1O1lIOOIlO0l01IIIIII,IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII,IO0010l0I011lIOIOOl1O1l101lllIIIII,IOOOOOl1OOO010IO00O0IO0Il10O1IIIII
,IO1IOI00OI0I10OO1l0I0l1l010llIIIII);IO10I111l1OOlIO0IlI1I00llll0lIIIII:=TRUE;END IF;WHEN OTHERS=>NULL;END CASE;IF IO10I111l1OOlIO0IlI1I00llll0lIIIII THEN IOOl0O0Il1Il00ll0l0l110I1OIllIIIII:=IIOO10OO0IlIl1l0II1O1lOIOI0IlIIIII;IIO0lO00IO0IO01O001OIOlll11OlIIIII:=
IO0010l0I011lIOIOOl1O1l101lllIIIII;II000llI0IIOIlO0OO01I11I01000IIIII:=IOOOOOl1OOO010IO00O0IO0Il10O1IIIII;II1IIlIllI0l0O110Il0OlIII1OOOIIIII:=IO1IOI00OI0I10OO1l0I0l1l010llIIIII;IIO0ll0III00OIOOI1I1OI1lIlO1OIIIII:=IOllIl0O0Ollll0IOlI011lI01Il1IIIII;ELSE IOOl0O0Il1Il00ll0l0l110I1OIllIIIII:=(OTHERS=>'X');
IIO0lO00IO0IO01O001OIOlll11OlIIIII:='X';II000llI0IIOIlO0OO01I11I01000IIIII:='X';II1IIlIllI0l0O110Il0OlIII1OOOIIIII:='X';IIO0ll0III00OIOOI1I1OI1lIlO1OIIIII:='X';END IF;END;CONSTANT IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII:GENERICS_TYPE:=
FLOATING_POINT_V6_0_CHECK_GENERICS(C_XDEVICEFAMILY=>C_XDEVICEFAMILY,C_HAS_ADD=>C_HAS_ADD,C_HAS_SUBTRACT=>C_HAS_SUBTRACT,
C_HAS_MULTIPLY=>C_HAS_MULTIPLY,C_HAS_DIVIDE=>C_HAS_DIVIDE,C_HAS_SQRT=>C_HAS_SQRT,C_HAS_COMPARE=>C_HAS_COMPARE,C_HAS_FIX_TO_FLT=>
C_HAS_FIX_TO_FLT,C_HAS_FLT_TO_FIX=>C_HAS_FLT_TO_FIX,C_HAS_FLT_TO_FLT=>C_HAS_FLT_TO_FLT,C_HAS_RECIP=>C_HAS_RECIP,C_HAS_RECIP_SQRT=>
C_HAS_RECIP_SQRT,C_A_WIDTH=>C_A_WIDTH,C_A_FRACTION_WIDTH=>C_A_FRACTION_WIDTH,C_B_WIDTH=>C_B_WIDTH,C_B_FRACTION_WIDTH=>
C_B_FRACTION_WIDTH,C_RESULT_WIDTH=>C_RESULT_WIDTH,C_RESULT_FRACTION_WIDTH=>C_RESULT_FRACTION_WIDTH,C_COMPARE_OPERATION=>
C_COMPARE_OPERATION,C_LATENCY=>C_LATENCY,C_OPTIMIZATION=>C_OPTIMIZATION,C_MULT_USAGE=>C_MULT_USAGE,C_RATE=>C_RATE,C_HAS_UNDERFLOW=>
C_HAS_UNDERFLOW,C_HAS_OVERFLOW=>C_HAS_OVERFLOW,C_HAS_INVALID_OP=>C_HAS_INVALID_OP,C_HAS_DIVIDE_BY_ZERO=>C_HAS_DIVIDE_BY_ZERO,
C_HAS_ACLKEN=>C_HAS_ACLKEN,C_HAS_ARESETN=>C_HAS_ARESETN,C_THROTTLE_SCHEME=>C_THROTTLE_SCHEME,C_HAS_A_TUSER=>C_HAS_A_TUSER,
C_HAS_A_TLAST=>C_HAS_A_TLAST,C_HAS_B=>C_HAS_B,C_HAS_B_TUSER=>C_HAS_B_TUSER,C_HAS_B_TLAST=>C_HAS_B_TLAST,C_HAS_OPERATION=>
C_HAS_OPERATION,C_HAS_OPERATION_TUSER=>C_HAS_OPERATION_TUSER,C_HAS_OPERATION_TLAST=>C_HAS_OPERATION_TLAST,C_HAS_RESULT_TUSER=>
C_HAS_RESULT_TUSER,C_HAS_RESULT_TLAST=>C_HAS_RESULT_TLAST,C_TLAST_RESOLUTION=>C_TLAST_RESOLUTION,C_A_TDATA_WIDTH=>C_A_TDATA_WIDTH,
C_A_TUSER_WIDTH=>C_A_TUSER_WIDTH,C_B_TDATA_WIDTH=>C_B_TDATA_WIDTH,C_B_TUSER_WIDTH=>C_B_TUSER_WIDTH,C_OPERATION_TDATA_WIDTH=>
C_OPERATION_TDATA_WIDTH,C_OPERATION_TUSER_WIDTH=>C_OPERATION_TUSER_WIDTH,C_RESULT_TDATA_WIDTH=>C_RESULT_TDATA_WIDTH,
C_RESULT_TUSER_WIDTH=>C_RESULT_TUSER_WIDTH);CONSTANT IOllIl10l0Ol0OIIOI1110lI01IOOIIIII:STD_LOGIC_VECTOR(FLT_PT_OP_CODE_SLICE):=FLT_PT_GET_OP_CODE(
C_HAS_ADD=>C_HAS_ADD,C_HAS_SUBTRACT=>C_HAS_SUBTRACT,C_HAS_MULTIPLY=>C_HAS_MULTIPLY,C_HAS_DIVIDE=>C_HAS_DIVIDE,C_HAS_SQRT=>C_HAS_SQRT
,C_HAS_COMPARE=>C_HAS_COMPARE,C_HAS_FIX_TO_FLT=>C_HAS_FIX_TO_FLT,C_HAS_FLT_TO_FIX=>C_HAS_FLT_TO_FIX,C_HAS_FLT_TO_FLT=>
C_HAS_FLT_TO_FLT,C_HAS_RECIP=>C_HAS_RECIP,C_HAS_RECIP_SQRT=>C_HAS_RECIP_SQRT);CONSTANT IO1O1lll1OIO1100I0OI011OlO1I0IIIII:INTEGER:=FLT_PT_DELAY(FAMILY=>
C_XDEVICEFAMILY,OP_CODE=>IOllIl10l0Ol0OIIOI1110lI01IOOIIIII,A_WIDTH=>C_A_WIDTH,A_FRACTION_WIDTH=>C_A_FRACTION_WIDTH,B_WIDTH=>C_B_WIDTH,B_FRACTION_WIDTH=>
C_B_FRACTION_WIDTH,RESULT_WIDTH=>C_RESULT_WIDTH,RESULT_FRACTION_WIDTH=>C_RESULT_FRACTION_WIDTH,OPTIMIZATION=>C_OPTIMIZATION,
MULT_USAGE=>C_MULT_USAGE,RATE=>C_RATE,THROTTLE_SCHEME=>C_THROTTLE_SCHEME,HAS_ADD=>C_HAS_ADD,HAS_SUBTRACT=>C_HAS_SUBTRACT,
HAS_MULTIPLY=>C_HAS_MULTIPLY,HAS_DIVIDE=>C_HAS_DIVIDE,HAS_SQRT=>C_HAS_SQRT,HAS_COMPARE=>C_HAS_COMPARE,HAS_FLT_TO_FIX=>
C_HAS_FLT_TO_FIX,HAS_FIX_TO_FLT=>C_HAS_FIX_TO_FLT,HAS_FLT_TO_FLT=>C_HAS_FLT_TO_FLT,HAS_RECIP=>C_HAS_RECIP,HAS_RECIP_SQRT=>
C_HAS_RECIP_SQRT,REQUIRED=>C_LATENCY);FUNCTION IIOO1101O11lIlIIO1I0O1111OO1IOIIII(IOl11O00lO0I1Ol100IIOl11llI00IIIII:INTEGER)RETURN INTEGER IS CONSTANT
 IO01lI1I1I0I0l11101010Ol1ll11IIIII:INTEGER:=1;VARIABLE IIll1ll0lOl0OOl010OlI10lIII00IIIII:INTEGER:=0;BEGIN IF IOl11O00lO0I1Ol100IIOl11llI00IIIII/=CI_AND_TVALID_THROTTLE THEN IIll1ll0lOl0OOl010OlI10lIII00IIIII:=IIll1ll0lOl0OOl010OlI10lIII00IIIII+
IO01lI1I1I0I0l11101010Ol1ll11IIIII;END IF;RETURN IIll1ll0lOl0OOl010OlI10lIII00IIIII;END;CONSTANT IOl00O110IlO0Ol0l1111ll11011OIIIII:INTEGER:=IIOO1101O11lIlIIO1I0O1111OO1IOIIII(C_THROTTLE_SCHEME);
CONSTANT IIO01lOO1OlO00OlII0OIO1IOllI0IIIII:INTEGER:=2*BOOLEAN'pos(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE);CONSTANT IO11l1Ol0l11OOIlOOlO1O10OllllIIIII:INTEGER:=
IO1O1lll1OIO1100I0OI011OlO1I0IIIII-IOl00O110IlO0Ol0l1111ll11011OIIIII-IIO01lOO1OlO00OlII0OIO1IOllI0IIIII;SIGNAL IIl1O0l11lOOIOOIO1Il11O0O001IIIIII:STD_LOGIC:='0';SIGNAL IOlI011I01001IIOlOO00OIOOOlIIOIIII:STD_LOGIC:='1';SIGNAL
 IO01OOOO0lO0IOII11lI011OlOIl0IIIII:STD_LOGIC:='1';SIGNAL IO000OI1l1OlI0II10OO10O0101l0IIIII:STD_LOGIC:='0';SIGNAL IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII:STD_LOGIC:='0';SIGNAL II11111lIOOO1II00l01IIII0I11lIIIII:
STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II1OlO01OI01I0OIl1110OO11O0llIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_A_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IOO11OOOIII00O1I1lIIlII01OllIOIIII:STD_LOGIC:='0';SIGNAL IOOl0IOOO001O11l10OI01110l1O1IIIII:STD_LOGIC:='0';SIGNAL
 IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII:STD_LOGIC:='0';SIGNAL IO1IOIl1O1lII1IOI01IOI1O00IIOIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');
SIGNAL IIIOl1OlIOIOOOOO001I11lOI0O11IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II1OlI1ll1lI11OOl1llOI00O0lI1IIIII:STD_LOGIC:=
'0';SIGNAL IIIOlI1lOIIlI01l1I0IO1I010O10IIIII:STD_LOGIC:='0';SIGNAL IOOl010OO0lO0111O00l0Il1I1O1OIIIII:STD_LOGIC:='0';SIGNAL IOl01I0lI0II1l0l110IO011II0l1IIIII
:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IIO1I1O01lO0lOlI1lIl00O0Ol000IIIII:STD_LOGIC_VECTOR(
IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IO1l10OOlIlI011IIll1lI01I01OIIIIII:STD_LOGIC:='0';SIGNAL
 IIO00110IlIOl01O1I0O10100O111IIIII:STD_LOGIC:='0';SIGNAL II11O1O1I11O1l1OOlOll0O11I10IOIIII:STD_LOGIC:='0';SIGNAL IIO00110lO0OI1OOI01011ll0II0IOIIII:STD_LOGIC_VECTOR(
IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II001O10OO10OI0l00lOI0OlOI0IOIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_RESULT_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IOlOI0l01llI0OI011lO0010II101IIIII:STD_LOGIC:='0';SIGNAL IIOl0O00I1I01O00O1OlIO10I1l1IOIIII:STD_LOGIC_VECTOR(
IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IIOO1OlOIIIOIllOOOO1l1lI0OI0OIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_TUSER_WIDTH-1 DOWNTO 0):=(
OTHERS=>'0');SIGNAL II100001IOIO11OlIIlI0l1O1I1lIOIIII:STD_LOGIC:='0';SIGNAL IOllIll0010111OOOll10OO1l1OOlIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>
'0');SIGNAL IOlllllOII10I1OIII11111Oll010IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII:STD_LOGIC:='0';
SIGNAL IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IIIl0llII1l1II0llIOI1Ol00000OIIIII
:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL IIlOlO111l01IlO000Ol10Ol0O1I0IIIII:STD_LOGIC:='0';SIGNAL
 IOIIlOI0II0Ol11I1O11I10IOI111IIIII:STD_LOGIC:='0';SIGNAL IIIOOlIIlOO00lO1l11lI00O00OI1IIIII:STD_LOGIC:='0';SIGNAL IOOOOI11I0llOOl00OIII01l11I1IIIIII:STD_LOGIC:='1';SIGNAL IIll0l11IOll1011I1110l0lI1000IIIII:STD_LOGIC:='0';SIGNAL
 II1OOII1l0IOOOl0Oll1O0IIOO10OIIIII:STD_LOGIC:='0';SIGNAL IOIO10OIll1O1lO011I0OOl1I1OOIOIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TDATA_WIDTH-1 DOWNTO 0):=(OTHERS
=>'0');SIGNAL IO1IOI1Ol01O0I0llO1l0O010ll00IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TUSER_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');SIGNAL
 IOllOI0l1OI1IIO1II1l11IOll1l1IIIII:STD_LOGIC:='0';CONSTANT IO10OI11lI1I1Il0OI0l1IlI11Ol1IIIII:INTEGER:=1;CONSTANT IO1I1lI01ll001l0Il1lIll11O0O0IIIII:INTEGER:=IIO00110lO0OI1OOI01011ll0II0IOIIII'length
+II001O10OO10OI0l00lOI0OlOI0IOIIIII'length+IO10OI11lI1I1Il0OI0l1IlI11Ol1IIIII;SIGNAL IOOO0lIIO0Ol1Il10OI0lOl00IOl1IIIII:STD_LOGIC:='0';SIGNAL IOOO1IOOOIOIlO0Ol0l0O1OlI11I0IIIII,IOlOlIllOO00O1O1101001I11IlIlIIIII:STD_LOGIC_VECTOR(
IO1I1lI01ll001l0Il1lIll11O0O0IIIII-1 DOWNTO 0):=(OTHERS=>'0');PROCEDURE IO1IlO1O0l1llOOlOlIOlIIOI00I1IIIII(CONSTANT IO10IO10lOIOlO0l10OOOOII0O0l0IIIII:IN INTEGER;CONSTANT IOOl0Ol10Il101010O10lO0OOOIOIIIIII:IN BOOLEAN;
CONSTANT IOI1lOI11II111011ll10IO1IIOlIOIIII:IN BOOLEAN;II0I0OI01O11l100I1IOOOlO0I00OIIIII:IN STD_LOGIC_VECTOR;IIII00I11l1l0lO1IO11OI101O010IIIII:IN STD_LOGIC_VECTOR;IOlOI11lI11001lOIlI1lII0I0IIIOIIII:IN STD_LOGIC;SIGNAL III1Il1IOl0001I10lO1llO0l01O1IIIII:OUT
 STD_LOGIC_VECTOR)IS VARIABLE IIlO1ll1100I100OI01OIlOll0O1IOIIII:STD_LOGIC_VECTOR(IO10IO10lOIOlO0l10OOOOII0O0l0IIIII-1 DOWNTO 0);VARIABLE II1llOIlIO01IIlOIOIO10111l010IIIII:INTEGER:=0;BEGIN IIlO1ll1100I100OI01OIlOll0O1IOIIII(II0I0OI01O11l100I1IOOOlO0I00OIIIII'high
 DOWNTO 0):=II0I0OI01O11l100I1IOOOlO0I00OIIIII;II1llOIlIO01IIlOIOIO10111l010IIIII:=II0I0OI01O11l100I1IOOOlO0I00OIIIII'length;IF IOOl0Ol10Il101010O10lO0OOOIOIIIIII THEN IIlO1ll1100I100OI01OIlOll0O1IOIIII(IIII00I11l1l0lO1IO11OI101O010IIIII'high+II1llOIlIO01IIlOIOIO10111l010IIIII DOWNTO II1llOIlIO01IIlOIOIO10111l010IIIII):=IIII00I11l1l0lO1IO11OI101O010IIIII;II1llOIlIO01IIlOIOIO10111l010IIIII:=II1llOIlIO01IIlOIOIO10111l010IIIII+IIII00I11l1l0lO1IO11OI101O010IIIII'length;END IF;IF
 IOI1lOI11II111011ll10IO1IIOlIOIIII THEN IIlO1ll1100I100OI01OIlOll0O1IOIIII(II1llOIlIO01IIlOIOIO10111l010IIIII):=IOlOI11lI11001lOIlI1lII0I0IIIOIIII;END IF;III1Il1IOl0001I10lO1llO0l01O1IIIII<=IIlO1ll1100I100OI01OIlOll0O1IOIIII;END;PROCEDURE IOO0O1IlI1O11O01O111010Ol10lOIIIII(CONSTANT IO10I1lIll0I0lO0IO1lOIIOIO0lIIIIII:IN INTEGER
;CONSTANT IO0O01O0IO0lOO1l001O10O100100IIIII:IN BOOLEAN;CONSTANT IIlOIl1000I0llI0llOIIllO11lOOIIIII:IN BOOLEAN;SIGNAL IIOI000I11lOl0OO1l01Oll1IlO1lIIIII:IN STD_LOGIC_VECTOR;SIGNAL IIOOI00000OO00O10l1lOIIIOl1lIOIIII:OUT
 STD_LOGIC_VECTOR;SIGNAL IO10O0OI111O0III0OI0Ol0I0llOOIIIII:OUT STD_LOGIC_VECTOR;SIGNAL IOOllO1OO0IlII00llll11I1IIO1IIIIII:OUT STD_LOGIC)IS VARIABLE IO0IIO01IIOIlOllO110l0l0010OlIIIII:INTEGER:=0;BEGIN IIOOI00000OO00O10l1lOIIIOl1lIOIIII<=IIOI000I11lOl0OO1l01Oll1IlO1lIIIII
(IIOOI00000OO00O10l1lOIIIOl1lIOIIII'high DOWNTO 0);IO0IIO01IIOIlOllO110l0l0010OlIIIII:=IIOOI00000OO00O10l1lOIIIOl1lIOIIII'length;IF IO0O01O0IO0lOO1l001O10O100100IIIII THEN IO10O0OI111O0III0OI0Ol0I0llOOIIIII<=IIOI000I11lOl0OO1l01Oll1IlO1lIIIII(IO10O0OI111O0III0OI0Ol0I0llOOIIIII'high+IO0IIO01IIOIlOllO110l0l0010OlIIIII DOWNTO IO0IIO01IIOIlOllO110l0l0010OlIIIII);IO0IIO01IIOIlOllO110l0l0010OlIIIII:=IO0IIO01IIOIlOllO110l0l0010OlIIIII+IO10O0OI111O0III0OI0Ol0I0llOOIIIII'length;END
 IF;IF IIlOIl1000I0llI0llOIIllO11lOOIIIII THEN IOOllO1OO0IlII00llll11I1IIO1IIIIII<=IIOI000I11lOl0OO1l01Oll1IlO1lIIIII(IO0IIO01IIOIlOllO110l0l0010OlIIIII);END IF;END;SIGNAL IOlII01I0000OII0I1OIO0I0OIO10IIIII:STD_LOGIC_VECTOR(IIO00110lO0OI1OOI01011ll0II0IOIIII'range
):=(OTHERS=>'0');SIGNAL IOllOlO0II0IIOlOOIOlI1l0OOIOIOIIII:STD_LOGIC_VECTOR(II001O10OO10OI0l00lOI0OlOI0IOIIIII'range):=(OTHERS=>'0');SIGNAL
 IO1II000OlOO0lOO1O0OI0lI1Il1OIIIII:STD_LOGIC:='0';SIGNAL IO0l0110O110I1I0O01I000ll11O1IIIII:STD_LOGIC:='0';SIGNAL II01ll1IOIO0110II0O0OlOIO110lIIIII:STD_LOGIC:='0';BEGIN
 IIl1O0l11lOOIOOIO1Il11O0O001IIIIII<=ACLK;IOlI011I01001IIOlOO00OIOOOlIIOIIII<=ACLKEN WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_ACLKEN=1 ELSE '1';IO01OOOO0lO0IOII11lI011OlOIl0IIIII<=ARESETN WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_ARESETN=1 ELSE '1'
;IO000OI1l1OlI0II10OO10O0101l0IIIII<=S_AXIS_A_TVALID;II11111lIOOO1II00l01IIII0I11lIIIII<=S_AXIS_A_TDATA;II1OlO01OI01I0OIl1110OO11O0llIIIII<=S_AXIS_A_TUSER WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TUSER
=1 ELSE(OTHERS=>'0');IOO11OOOIII00O1I1lIIlII01OllIOIIII<=S_AXIS_A_TLAST WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TLAST=1 ELSE '0';IOOl0IOOO001O11l10OI01110l1O1IIIII<=S_AXIS_B_TVALID
 WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B=1 ELSE '1';IO1IOIl1O1lII1IOI01IOI1O00IIOIIIII<=S_AXIS_B_TDATA WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B=1 ELSE(OTHERS=>'0');IIIOl1OlIOIOOOOO001I11lOI0O11IIIII
<=S_AXIS_B_TUSER WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TUSER=1 ELSE(OTHERS=>'0');II1OlI1ll1lI11OOl1llOI00O0lI1IIIII<=S_AXIS_B_TLAST WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TLAST
=1 ELSE '0';IIIOlI1lOIIlI01l1I0IO1I010O10IIIII<=S_AXIS_OPERATION_TVALID WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION=1 ELSE '1';IOl01I0lI0II1l0l110IO011II0l1IIIII
<=S_AXIS_OPERATION_TDATA WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION=1 ELSE(OTHERS=>'0');IIO1I1O01lO0lOlI1lIl00O0Ol000IIIII<=S_AXIS_OPERATION_TUSER WHEN
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION_TUSER=1 ELSE(OTHERS=>'0');IO1l10OOlIlI011IIll1lI01I01OIIIIII<=S_AXIS_OPERATION_TLAST WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_OPERATION_TLAST=1 ELSE '0';II11O1O1I11O1l1OOlOll0O11I10IOIIII<=M_AXIS_RESULT_TREADY WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE OR
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_CE_THROTTLE)ELSE '1';REG_SCLR:PROCESS(ACLK)BEGIN IF RISING_EDGE(ACLK)THEN IIll0l11IOll1011I1110l0lI1000IIIII<=NOT IO01OOOO0lO0IOII11lI011OlOIl0IIIII;END
 IF;END PROCESS;AND_TVALIDS_CTRL:IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE GENERATE SIGNAL IIOI0110I1IOI00OOl01IO0I0O0IIOIIII:INTEGER:=0;
BEGIN IIOl0O00I1I01O00O1OlIO10I1l1IOIIII<=II11111lIOOO1II00l01IIII0I11lIIIII;IIOO1OlOIIIOIllOOOO1l1lI0OI0OIIIII<=II1OlO01OI01I0OIl1110OO11O0llIIIII;II100001IOIO11OlIIlI0l1O1I1lIOIIII<=IOO11OOOIII00O1I1lIIlII01OllIOIIII;IOllIll0010111OOOll10OO1l1OOlIIIII<=IO1IOIl1O1lII1IOI01IOI1O00IIOIIIII;IOlllllOII10I1OIII11111Oll010IIIII
<=IIIOl1OlIOIOOOOO001I11lOI0O11IIIII;II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII<=II1OlI1ll1lI11OOl1llOI00O0lI1IIIII;IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII<=IOl01I0lI0II1l0l110IO011II0l1IIIII;IIIl0llII1l1II0llIOI1Ol00000OIIIII<=
IIO1I1O01lO0lOlI1lIl00O0Ol000IIIII;IIlOlO111l01IlO000Ol10Ol0O1I0IIIII<=IO1l10OOlIlI011IIll1lI01I01OIIIIII;IOIIlOI0II0Ol11I1O11I10IOI111IIIII<=IO000OI1l1OlI0II10OO10O0101l0IIIII AND IOOl0IOOO001O11l10OI01110l1O1IIIII AND
 IIIOlI1lOIIlI01l1I0IO1I010O10IIIII;IIIOOlIIlOO00lO1l11lI00O00OI1IIIII<='0';LATENCY_GT_ZERO:IF C_LATENCY>0 GENERATE RATE_COUNTER:PROCESS(ACLK)BEGIN IF RISING_EDGE
(ACLK)THEN IF IIll0l11IOll1011I1110l0lI1000IIIII='1'THEN IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1 THEN IOOOOI11I0llOOl00OIII01l11I1IIIIII<='0';END IF;IIOI0110I1IOI00OOl01IO0I0O0IIOIIII<=0;IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII<='0';
IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII<='0';IOOl010OO0lO0111O00l0Il1I1O1OIIIII<='0';ELSIF IOlI011I01001IIOlOO00OIOOOlIIOIIII='1'THEN IF IIOI0110I1IOI00OOl01IO0I0O0IIOIIII=0 THEN IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII<='1';
IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII<='1';IOOl010OO0lO0111O00l0Il1I1O1OIIIII<='1';ELSE IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII<='0';IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII<='0';IOOl010OO0lO0111O00l0Il1I1O1OIIIII
<='0';END IF;IF IIOI0110I1IOI00OOl01IO0I0O0IIOIIII=0 THEN IIOI0110I1IOI00OOl01IO0I0O0IIOIIII<=IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE-1;ELSE IIOI0110I1IOI00OOl01IO0I0O0IIOIIII<=IIOI0110I1IOI00OOl01IO0I0O0IIOIIII-1;END IF;IF
 IIOI0110I1IOI00OOl01IO0I0O0IIOIIII=0 THEN IOOOOI11I0llOOl00OIII01l11I1IIIIII<='1';ELSE IOOOOI11I0llOOl00OIII01l11I1IIIIII<='0';END IF;END IF;END IF;END PROCESS;END GENERATE;LATENCY_ZERO:IF C_LATENCY=0
 GENERATE IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII<='1';IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII<='1';IOOl010OO0lO0111O00l0Il1I1O1OIIIII<='1';IOOOOI11I0llOOl00OIII01l11I1IIIIII<='1';END GENERATE;END GENERATE;
AXI_CTRL:IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME/=CI_AND_TVALID_THROTTLE GENERATE CONSTANT IO0lO0Il1IlIllI1O0OI1l0lO10I0IIIII:BOOLEAN:=NOT(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_THROTTLE_SCHEME=CI_GEN_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE=1);SIGNAL IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII:INTEGER:=0;SIGNAL IIIlOl1O101100O0OOl00l1l1OlOOIIIII:STD_LOGIC:='0';
SIGNAL IOllI11l100l00I101O100Il100IOOIIII:STD_LOGIC;SIGNAL II00O0lIIO0IlIIII10l010I1001OIIIII:STD_LOGIC_VECTOR(C_A_TDATA_WIDTH-1 DOWNTO 0);SIGNAL IIIIlO11IO11lI1OII0l0IO0IlI1lIIIII:STD_LOGIC_VECTOR(
C_A_TUSER_WIDTH-1 DOWNTO 0);SIGNAL II1II1O0OOI00111l1Il1O10l1Il0IIIII:STD_LOGIC;SIGNAL IIIO0O11100l00l110OlOOIII00lIOIIII:STD_LOGIC_VECTOR(C_B_TDATA_WIDTH-1 DOWNTO 0);SIGNAL
 II1I0Il1010l11l00I10lII0l0l10IIIII:STD_LOGIC_VECTOR(C_B_TUSER_WIDTH-1 DOWNTO 0);SIGNAL IOI11I1I0I1IOI0llIO11101IOlOIOIIII:STD_LOGIC;SIGNAL IOOI01O1OlO11OOOlOIll1OI101IlIIIII:
STD_LOGIC_VECTOR(C_OPERATION_TDATA_WIDTH-1 DOWNTO 0);SIGNAL II1l0Ol0O0lO101IO110011O11IOOIIIII:STD_LOGIC_VECTOR(C_OPERATION_TUSER_WIDTH-1 DOWNTO 0
);SIGNAL IOI11Oll1O010II0IlIOI0IO01IIlIIIII:STD_LOGIC;BEGIN I_SYNC:AXI_SLAVE_3TO1_V1_1 GENERIC MAP(C_A_TDATA_WIDTH=>C_A_TDATA_WIDTH,C_HAS_A_TUSER
=>C_HAS_A_TUSER=1,C_A_TUSER_WIDTH=>C_A_TUSER_WIDTH,C_HAS_A_TLAST=>C_HAS_A_TLAST=1,C_B_TDATA_WIDTH=>C_B_TDATA_WIDTH,C_HAS_B_TUSER=>
C_HAS_B_TUSER=1,C_B_TUSER_WIDTH=>C_B_TUSER_WIDTH,C_HAS_B_TLAST=>C_HAS_B_TLAST=1,C_C_TDATA_WIDTH=>C_OPERATION_TDATA_WIDTH,
C_HAS_C_TUSER=>C_HAS_OPERATION_TUSER=1,C_C_TUSER_WIDTH=>C_OPERATION_TUSER_WIDTH,C_HAS_C_TLAST=>C_HAS_OPERATION_TLAST=1,
C_HAS_Z_TREADY=>IO0lO0Il1IlIllI1O0OI1l0lO10I0IIIII)PORT MAP(ACLK,IOlI011I01001IIOlOO00OIOOOlIIOIIII,IIll0l11IOll1011I1110l0lI1000IIIII,IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII,IO000OI1l1OlI0II10OO10O0101l0IIIII,S_AXIS_A_TDATA,S_AXIS_A_TUSER,
S_AXIS_A_TLAST,IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII,IOOl0IOOO001O11l10OI01110l1O1IIIII,S_AXIS_B_TDATA,S_AXIS_B_TUSER,S_AXIS_B_TLAST,IOOl010OO0lO0111O00l0Il1I1O1OIIIII,
IIIOlI1lOIIlI01l1I0IO1I010O10IIIII,S_AXIS_OPERATION_TDATA,S_AXIS_OPERATION_TUSER,S_AXIS_OPERATION_TLAST,IIIlOl1O101100O0OOl00l1l1OlOOIIIII,IOllI11l100l00I101O100Il100IOOIIII,II00O0lIIO0IlIIII10l010I1001OIIIII
,IIIIlO11IO11lI1OII0l0IO0IlI1lIIIII,II1II1O0OOI00111l1Il1O10l1Il0IIIII,IIIO0O11100l00l110OlOOIII00lIOIIII,II1I0Il1010l11l00I10lII0l0l10IIIII,IOI11I1I0I1IOI0llIO11101IOlOIOIIII,IOOI01O1OlO11OOOlOIll1OI101IlIIIII,II1l0Ol0O0lO101IO110011O11IOOIIIII,IOI11Oll1O010II0IlIOI0IO01IIlIIIII);
IOIIlOI0II0Ol11I1O11I10IOI111IIIII<=IOllI11l100l00I101O100Il100IOOIIII;IIOl0O00I1I01O00O1OlIO10I1l1IOIIII<=II00O0lIIO0IlIIII10l010I1001OIIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_TDATA_WIDTH-1 DOWNTO 0);IIOO1OlOIIIOIllOOOO1l1lI0OI0OIIIII<=IIIIlO11IO11lI1OII0l0IO0IlI1lIIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_A_TUSER_WIDTH-1 DOWNTO 0)WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TUSER=1 ELSE(OTHERS=>'0');II100001IOIO11OlIIlI0l1O1I1lIOIIII<=II1II1O0OOI00111l1Il1O10l1Il0IIIII WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_A_TLAST=1 ELSE '0';IOllIll0010111OOOll10OO1l1OOlIIIII<=IIIO0O11100l00l110OlOOIII00lIOIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TDATA_WIDTH-1 DOWNTO 0);IOlllllOII10I1OIII11111Oll010IIIII<=II1I0Il1010l11l00I10lII0l0l10IIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_B_TUSER_WIDTH-1 DOWNTO 0)WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TUSER=1 ELSE(OTHERS=>'0');II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII<=IOI11I1I0I1IOI0llIO11101IOlOIOIIII WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_B_TLAST=1 ELSE '0';IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII<=IOOI01O1OlO11OOOlOIll1OI101IlIIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TDATA_WIDTH-1 DOWNTO 0);IIIl0llII1l1II0llIOI1Ol00000OIIIII
<=II1l0Ol0O0lO101IO110011O11IOOIIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TUSER_WIDTH-1 DOWNTO 0)WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION_TUSER=1 ELSE(OTHERS=>'0');
IIlOlO111l01IlO000Ol10Ol0O1I0IIIII<=IOI11Oll1O010II0IlIOI0IO01IIlIIIII WHEN IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION_TLAST=1 ELSE '0';RATE_COUNTER:PROCESS(ACLK)BEGIN IF
 RISING_EDGE(ACLK)THEN IF IIll0l11IOll1011I1110l0lI1000IIIII='1'THEN IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII<=0;ELSIF IOlI011I01001IIOlOO00OIOOOlIIOIIII='1'AND(IIIOOlIIlOO00lO1l11lI00O00OI1IIIII='0'OR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=
CI_RFD_THROTTLE AND IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII/=0))THEN IF IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII=0 THEN IF IOOOOI11I0llOOl00OIII01l11I1IIIIII='1'THEN IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII<=IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE-1;END IF
;ELSE IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII<=IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII-1;END IF;END IF;END IF;END PROCESS;IIIOOlIIlOO00lO1l11lI00O00OI1IIIII<='0'WHEN IIll0l11IOll1011I1110l0lI1000IIIII='1'ELSE IIO00110IlIOl01O1I0O10100O111IIIII
 AND NOT II11O1O1I11O1l1OOlOll0O11I10IOIIII;IIIlOl1O101100O0OOl00l1l1OlOOIIIII<=NOT IIIOOlIIlOO00lO1l11lI00O00OI1IIIII WHEN IOIlOl1I0I0OOI11lll0I0I01OI0OIIIII=0 ELSE '0';IOOOOI11I0llOOl00OIII01l11I1IIIIII<=IIIlOl1O101100O0OOl00l1l1OlOOIIIII AND IOIIlOI0II0Ol11I1O11I10IOI111IIIII;END
 GENERATE;CALC_RESULTS:PROCESS(IIIOOlIIlOO00lO1l11lI00O00OI1IIIII,IOOOOI11I0llOOl00OIII01l11I1IIIIII,IOIIlOI0II0Ol11I1O11I10IOI111IIIII,IIOl0O00I1I01O00O1OlIO10I1l1IOIIII,IOllIll0010111OOOll10OO1l1OOlIIIII,IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII,IIOO1OlOIIIOIllOOOO1l1lI0OI0OIIIII,IOlllllOII10I1OIII11111Oll010IIIII,
IIIl0llII1l1II0llIOI1Ol00000OIIIII,II100001IOIO11OlIIlI0l1O1I1lIOIIII,II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII,IIlOlO111l01IlO000Ol10Ol0O1I0IIIII)VARIABLE IIOIl1llO0OlI1l1llI1I0l11O1I0IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_WIDTH-1 DOWNTO 0):=(OTHERS
=>'0');VARIABLE IIO0Ol01I0lO11ll11O10OllOO001IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE IIIO1llOlO1II10II1O0llOIIOl1IIIIII:STD_LOGIC_VECTOR(
FLT_PT_OPERATION_WIDTH-1 DOWNTO 0):=(OTHERS=>'0');VARIABLE II0IOO0OI11010l0O1l1010IllO01IIIII:STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_WIDTH-1 DOWNTO 0):=(
OTHERS=>'0');VARIABLE II00OI01lllI1I1I1I0IIllOllIlIOIIII:STD_LOGIC:='0';VARIABLE IOO00OI0Il0O000lIlOOIllII1OOIIIIII:STD_LOGIC:='0';VARIABLE IIII1llI1I11lOI00IOOOIOl1OO0IIIIII:STD_LOGIC:='0'
;VARIABLE IIIllllI01O1110OO1l0I1lIII1O0IIIII:STD_LOGIC:='0';VARIABLE IOIOOl01l10O1llI1l00I01O1llIIIIIII:INTEGER:=0;BEGIN IF IIIOOlIIlOO00lO1l11lI00O00OI1IIIII='0'THEN II1OOII1l0IOOOl0Oll1O0IIOO10OIIIII<=
IOOOOI11I0llOOl00OIII01l11I1IIIIII AND IOIIlOI0II0Ol11I1O11I10IOI111IIIII;END IF;IF IOOOOI11I0llOOl00OIII01l11I1IIIIII='1'THEN IIOIl1llO0OlI1l1llI1I0l11O1I0IIIII:=IIOl0O00I1I01O00O1OlIO10I1l1IOIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_WIDTH-1 DOWNTO 0);IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B=1 THEN IIO0Ol01I0lO11ll11O10OllOO001IIIII:=
IOllIll0010111OOOll10OO1l1OOlIIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_WIDTH-1 DOWNTO 0);ELSE IIO0Ol01I0lO11ll11O10OllOO001IIIII:=(OTHERS=>'0');END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION=1 THEN IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_COMPARE=1 THEN IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_OP_CODE_SLICE):=FLT_PT_COMPARE_OP_CODE_SLV;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_COMPARE_OPERATION=
FLT_PT_PROGRAMMABLE THEN IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_COMPARE_OPERATION_SLICE):=FLT_PT_GET_COMPARE_OP(IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII(FLT_PT_OPERATION_WIDTH
-1 DOWNTO 0));ELSE IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_COMPARE_OPERATION_SLICE):=CONV_INT_TO_SLV_3(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_COMPARE_OPERATION,3);END IF;ELSIF
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_ADD=1 AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_SUBTRACT=1 THEN IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_OP_CODE_SLICE):=FLT_PT_ADD_OP_CODE_SLV;IIIO1llOlO1II10II1O0llOIIOl1IIIIII(0)
:=FLT_PT_GET_ADDSUB_OP(IOO001OIO1O1lIOO0OlOOOIO0O1OlIIIII(FLT_PT_OPERATION_WIDTH-1 DOWNTO 0));IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_COMPARE_OPERATION_SLICE):=(OTHERS=>
'0');ELSE REPORT"ERROR: floating_point_v6_0 behavioral model: unknown operators when OPERATION channel present"SEVERITY ERROR;END IF
;ELSE IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_OP_CODE_SLICE):=IOllIl10l0Ol0OIIOI1110lI01IOOIIIII;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_COMPARE=1 THEN IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_COMPARE_OPERATION_SLICE):=
CONV_INT_TO_SLV_3(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_COMPARE_OPERATION,3);ELSE IIIO1llOlO1II10II1O0llOIIOl1IIIIII(FLT_PT_COMPARE_OPERATION_SLICE):=(OTHERS=>'0');END IF;END IF;
II11l0O1IO1OOI000IIO11I1Oll1IIIIII(IOO011IOl1001I1O1lIOOIlO0l01IIIIII=>IIOIl1llO0OlI1l1llI1I0l11O1I0IIIII,IOIOIOOII1OO1I00OlOl1IIOll1OlIIIII=>IIO0Ol01I0lO11ll11O10OllOO001IIIII,IOlOII1IIOlI01OI0IOOIllI0I1IOIIIII=>IIIO1llOlO1II10II1O0llOIIOl1IIIIII,IOOl0O0Il1Il00ll0l0l110I1OIllIIIII=>II0IOO0OI11010l0O1l1010IllO01IIIII,IIO0lO00IO0IO01O001OIOlll11OlIIIII=>II00OI01lllI1I1I1I0IIllOllIlIOIIII,II000llI0IIOIlO0OO01I11I01000IIIII=>IOO00OI0Il0O000lIlOOIllII1OOIIIIII,II1IIlIllI0l0O110Il0OlIII1OOOIIIII=>
IIII1llI1I11lOI00IOOOIOl1OO0IIIIII,IIO0ll0III00OIOOI1I1OI1lIlO1OIIIII=>IIIllllI01O1110OO1l0I1lIII1O0IIIII);IOIO10OIll1O1lO011I0OOl1I1OOIOIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_WIDTH-1 DOWNTO 0)<=II0IOO0OI11010l0O1l1010IllO01IIIII;IF
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_COMPARE=1 THEN IOIO10OIll1O1lO011I0OOl1I1OOIOIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TDATA_WIDTH-1 DOWNTO IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_WIDTH)<=(OTHERS
=>'0');ELSE IOIO10OIll1O1lO011I0OOl1I1OOIOIIII(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TDATA_WIDTH-1 DOWNTO IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_WIDTH)<=(OTHERS=>II0IOO0OI11010l0O1l1010IllO01IIIII(
II0IOO0OI11010l0O1l1010IllO01IIIII'left));END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TUSER=1 THEN IOIOOl01l10O1llI1l00I01O1llIIIIIII:=0;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_UNDERFLOW=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IIII1llI1I11lOI00IOOOIOl1OO0IIIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+1;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OVERFLOW=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IOO00OI0Il0O000lIlOOIllII1OOIIIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+1;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_INVALID_OP=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=II00OI01lllI1I1I1I0IIllOllIlIOIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+1;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_DIVIDE_BY_ZERO=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IIIllllI01O1110OO1l0I1lIII1O0IIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+1;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TUSER=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII+IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_A_TUSER_WIDTH-1 DOWNTO IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IIOO1OlOIIIOIllOOOO1l1lI0OI0OIIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_A_TUSER_WIDTH;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TUSER=1 THEN IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII+IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TUSER_WIDTH-1 DOWNTO
 IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IOlllllOII10I1OIII11111Oll010IIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_B_TUSER_WIDTH;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION_TUSER=1 THEN
 IO1IOI1Ol01O0I0llO1l0O010ll00IIIII(IOIOOl01l10O1llI1l00I01O1llIIIIIII+IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TUSER_WIDTH-1 DOWNTO IOIOOl01l10O1llI1l00I01O1llIIIIIII)<=IIIl0llII1l1II0llIOI1Ol00000OIIIII;IOIOOl01l10O1llI1l00I01O1llIIIIIII:=IOIOOl01l10O1llI1l00I01O1llIIIIIII+
IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_OPERATION_TUSER_WIDTH;END IF;ASSERT IOIOOl01l10O1llI1l00I01O1llIIIIIII=IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TUSER_WIDTH REPORT
"ERROR: floating_point_v6_0 behavioral model: Did not concatenate the correct number of bits "&
"when constructing m_axis_result_tuser: expected "&INTEGER'image(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TUSER_WIDTH)&", actual "&INTEGER'image(
IOIOOl01l10O1llI1l00I01O1llIIIIIII)SEVERITY ERROR;END IF;IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TLAST=1 THEN CASE IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_TLAST_RESOLUTION IS WHEN CI_TLAST_PASS_A
=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII<=II100001IOIO11OlIIlI0l1O1I1lIOIIII;WHEN CI_TLAST_PASS_B=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII<=II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII;WHEN CI_TLAST_PASS_C=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII<=
IIlOlO111l01IlO000Ol10Ol0O1I0IIIII;WHEN CI_TLAST_OR_ALL=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII<=((II100001IOIO11OlIIlI0l1O1I1lIOIIII AND CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TLAST=1))OR(
II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII AND CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TLAST=1))OR(IIlOlO111l01IlO000Ol10Ol0O1I0IIIII AND CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_OPERATION_TLAST=1)));WHEN CI_TLAST_AND_ALL=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII<=((II100001IOIO11OlIIlI0l1O1I1lIOIIII OR NOT CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_A_TLAST
=1))AND(II0lI1II01IlOIIOl1I1ll0I0I1IIIIIII OR NOT CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B_TLAST=1))AND(IIlOlO111l01IlO000Ol10Ol0O1I0IIIII OR NOT CONV_BOOL_TO_SL(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_OPERATION_TLAST=1)));WHEN OTHERS=>REPORT"ERROR: floating_point_v6_0 behavioral model: Unknown value of C_TLAST_RESOLUTION: "&
INTEGER'image(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_TLAST_RESOLUTION)SEVERITY ERROR;END CASE;END IF;END IF;END PROCESS;DELAY_0:IF IO11l1Ol0l11OOIlOOlO1O10OllllIIIII=0 GENERATE
 IO0l0110O110I1I0O01I000ll11O1IIIII<=II1OOII1l0IOOOl0Oll1O0IIOO10OIIIII;IOlII01I0000OII0I1OIO0I0OIO10IIIII<=IOIO10OIll1O1lO011I0OOl1I1OOIOIIII;IOllOlO0II0IIOlOOIOlI1l0OOIOIOIIII<=
IO1IOI1Ol01O0I0llO1l0O010ll00IIIII;IO1II000OlOO0lOO1O0OI0lI1Il1OIIIII<=IOllOI0l1OI1IIO1II1l11IOll1l1IIIII;IOOO0lIIO0Ol1Il10OI0lOl00IOl1IIIII<=IOOOOI11I0llOOl00OIII01l11I1IIIIII AND IOlI011I01001IIOlOO00OIOOOlIIOIIII;IO1IlO1O0l1llOOlOlIOlIIOI00I1IIIII(IO10IO10lOIOlO0l10OOOOII0O0l0IIIII=>
IO1I1lI01ll001l0Il1lIll11O0O0IIIII,IOOl0Ol10Il101010O10lO0OOOIOIIIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TUSER=1),IOI1lOI11II111011ll10IO1IIOlIOIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TLAST=1),II0I0OI01O11l100I1IOOOlO0I00OIIIII=>
IOIO10OIll1O1lO011I0OOl1I1OOIOIIII,IIII00I11l1l0lO1IO11OI101O010IIIII=>IO1IOI1Ol01O0I0llO1l0O010ll00IIIII,IOlOI11lI11001lOIlI1lII0I0IIIOIIII=>IOllOI0l1OI1IIO1II1l11IOll1l1IIIII,III1Il1IOl0001I10lO1llO0l01O1IIIII=>IOOO1IOOOIOIlO0Ol0l0O1OlI11I0IIIII);END GENERATE;DELAY_N:IF IO11l1Ol0l11OOIlOOlO1O10OllllIIIII/=0
 GENERATE MODEL:PROCESS(ACLK)TYPE IOO1l0lO1Il1l0OlOIOlO0OOllO1lIIIII IS ARRAY(NATURAL RANGE<>)OF STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TDATA_WIDTH-1
 DOWNTO 0);TYPE IIIllll0OIOl000lO1Il10OlI0OOlIIIII IS ARRAY(NATURAL RANGE<>)OF STD_LOGIC_VECTOR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RESULT_TUSER_WIDTH-1 DOWNTO 0);VARIABLE
 II01I1l01OOO10I00I000l0l0lI1IIIIII:STD_LOGIC_VECTOR(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII):=(OTHERS=>'0');VARIABLE II1O0lIl010OOll1OIO1IIOOlO1lIOIIII:IOO1l0lO1Il1l0OlOIOlO0OOllO1lIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII):=(OTHERS=>(OTHERS=>'0'));
VARIABLE IO00OlI1I01OOOOOIl100l0II0OIOIIIII:IIIllll0OIOl000lO1Il10OlI0OOlIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII):=(OTHERS=>(OTHERS=>'0'));VARIABLE II1111I0II10Ol0O01101I0O0000IIIIII:STD_LOGIC_VECTOR(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII):=(OTHERS
=>'0');VARIABLE II0O0O01lIOOlOl0IOllI1ll1O0I0IIIII:STD_LOGIC_VECTOR(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII):=(OTHERS=>'0');BEGIN IF RISING_EDGE(ACLK)THEN IF IIll0l11IOll1011I1110l0lI1000IIIII='1'THEN
 II01I1l01OOO10I00I000l0l0lI1IIIIII:=(OTHERS=>'0');IO0l0110O110I1I0O01I000ll11O1IIIII<='0';II0O0O01lIOOlOl0IOllI1ll1O0I0IIIII:=(OTHERS=>'0');II01ll1IOIO0110II0O0OlOIO110lIIIII<='0';ELSIF IOlI011I01001IIOlOO00OIOOOlIIOIIII='1'THEN
 II0O0O01lIOOlOl0IOllI1ll1O0I0IIIII:=IOOOOI11I0llOOl00OIII01l11I1IIIIII&II0O0O01lIOOlOl0IOllI1ll1O0I0IIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);II01ll1IOIO0110II0O0OlOIO110lIIIII<=II0O0O01lIOOlOl0IOllI1ll1O0I0IIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII);IF IIIOOlIIlOO00lO1l11lI00O00OI1IIIII='0'OR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_THROTTLE_SCHEME=CI_RFD_THROTTLE)THEN II01I1l01OOO10I00I000l0l0lI1IIIIII:=II1OOII1l0IOOOl0Oll1O0IIOO10OIIIII&II01I1l01OOO10I00I000l0l0lI1IIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);IO0l0110O110I1I0O01I000ll11O1IIIII<=
II01I1l01OOO10I00I000l0l0lI1IIIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII);END IF;END IF;IF(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE)THEN IF IOlI011I01001IIOlOO00OIOOOlIIOIIII='1'THEN II1O0lIl010OOll1OIO1IIOOlO1lIOIIII:=
IOIO10OIll1O1lO011I0OOl1I1OOIOIIII&II1O0lIl010OOll1OIO1IIOOlO1lIOIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);IO00OlI1I01OOOOOIl100l0II0OIOIIIII:=IO1IOI1Ol01O0I0llO1l0O010ll00IIIII&IO00OlI1I01OOOOOIl100l0II0OIOIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);II1111I0II10Ol0O01101I0O0000IIIIII:=
IOllOI0l1OI1IIO1II1l11IOll1l1IIIII&II1111I0II10Ol0O01101I0O0000IIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);IO1IlO1O0l1llOOlOlIOlIIOI00I1IIIII(IO10IO10lOIOlO0l10OOOOII0O0l0IIIII=>IO1I1lI01ll001l0Il1lIll11O0O0IIIII,IOOl0Ol10Il101010O10lO0OOOIOIIIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TUSER
=1),IOI1lOI11II111011ll10IO1IIOlIOIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TLAST=1),II0I0OI01O11l100I1IOOOlO0I00OIIIII=>II1O0lIl010OOll1OIO1IIOOlO1lIOIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII),IIII00I11l1l0lO1IO11OI101O010IIIII=>IO00OlI1I01OOOOOIl100l0II0OIOIIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII),IOlOI11lI11001lOIlI1lII0I0IIIOIIII=>II1111I0II10Ol0O01101I0O0000IIIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII),
III1Il1IOl0001I10lO1llO0l01O1IIIII=>IOOO1IOOOIOIlO0Ol0l0O1OlI11I0IIIII);END IF;ELSE IF IOlI011I01001IIOlOO00OIOOOlIIOIIII='1'THEN IF IIIOOlIIlOO00lO1l11lI00O00OI1IIIII='0'THEN II1O0lIl010OOll1OIO1IIOOlO1lIOIIII:=IOIO10OIll1O1lO011I0OOl1I1OOIOIIII&II1O0lIl010OOll1OIO1IIOOlO1lIOIIII(1 TO
 IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);IO00OlI1I01OOOOOIl100l0II0OIOIIIII:=IO1IOI1Ol01O0I0llO1l0O010ll00IIIII&IO00OlI1I01OOOOOIl100l0II0OIOIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);II1111I0II10Ol0O01101I0O0000IIIIII:=IOllOI0l1OI1IIO1II1l11IOll1l1IIIII&II1111I0II10Ol0O01101I0O0000IIIIII(1 TO IO11l1Ol0l11OOIlOOlO1O10OllllIIIII-1);
IOlII01I0000OII0I1OIO0I0OIO10IIIII<=II1O0lIl010OOll1OIO1IIOOlO1lIOIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII);IOllOlO0II0IIOlOOIOlI1l0OOIOIOIIII<=IO00OlI1I01OOOOOIl100l0II0OIOIIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII);IO1II000OlOO0lOO1O0OI0lI1Il1OIIIII<=
II1111I0II10Ol0O01101I0O0000IIIIII(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII);END IF;END IF;END IF;END IF;END PROCESS;IOOO0lIIO0Ol1Il10OI0lOl00IOl1IIIII<=II01ll1IOIO0110II0O0OlOIO110lIIIII AND IOlI011I01001IIOlOO00OIOOOlIIOIIII;END GENERATE;NO_OUTPUT_FIFO:IF
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME/=CI_RFD_THROTTLE GENERATE IIO00110lO0OI1OOI01011ll0II0IOIIII<=IOlII01I0000OII0I1OIO0I0OIO10IIIII;II001O10OO10OI0l00lOI0OlOI0IOIIIII<=
IOllOlO0II0IIOlOOIOlI1l0OOIOIOIIII;IOlOI0l01llI0OI011lO0010II101IIIII<=IO1II000OlOO0lOO1O0OI0lI1Il1OIIIII;IIO00110IlIOl01O1I0O10100O111IIIII<=IO0l0110O110I1I0O01I000ll11O1IIIII;END
 GENERATE;HAS_OUTPUT_FIFO:IF IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE GENERATE CONSTANT IIO01lO00lO0IllIOlllI11I0I1IIIIIII:INTEGER:=16;CONSTANT
 II1O0ll1Il100O1IIlOll0I00l1OOIIIII:INTEGER:=1;CONSTANT IIIO011I0OO0I0OIOl0llO11111OIOIIII:INTEGER:=FLT_PT_MAX(2**LOG2ROUNDUP(IO11l1Ol0l11OOIlOOlO1O10OllllIIIII+II1O0ll1Il100O1IIlOll0I00l1OOIIIII),IIO01lO00lO0IllIOlllI11I0I1IIIIIII);BEGIN
 OUTPUT_FIFO:GLB_IFX_MASTER_V1_1 GENERIC MAP(WIDTH=>IO1I1lI01ll001l0Il1lIll11O0O0IIIII,DEPTH=>IIIO011I0OO0I0OIOl0llO11111OIOIIII,AFULL_THRESH1=>1,AFULL_THRESH0=>1)
PORT MAP(ACLK=>ACLK,ACLKEN=>IOlI011I01001IIOlOO00OIOOOlIIOIIII,ARESET=>IIll0l11IOll1011I1110l0lI1000IIIII,WR_ENABLE=>IOOO0lIIO0Ol1Il10OI0lOl00IOl1IIIII,WR_DATA=>IOOO1IOOOIOIlO0Ol0l0O1OlI11I0IIIII,IFX_VALID=>IIO00110IlIOl01O1I0O10100O111IIIII,
IFX_READY=>M_AXIS_RESULT_TREADY,IFX_DATA=>IOlOlIllOO00O1O1101001I11IlIlIIIII,FULL=>OPEN,AFULL=>OPEN,NOT_FULL=>OPEN,NOT_AFULL=>OPEN,ADD=>OPEN);
IOO0O1IlI1O11O01O111010Ol10lOIIIII(IO10I1lIll0I0lO0IO1lOIIOIO0lIIIIII=>IO1I1lI01ll001l0Il1lIll11O0O0IIIII,IO0O01O0IO0lOO1l001O10O100100IIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TUSER=1),IIlOIl1000I0llI0llOIIllO11lOOIIIII=>(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_RESULT_TLAST=1),IIOI000I11lOl0OO1l01Oll1IlO1lIIIII=>IOlOlIllOO00O1O1101001I11IlIlIIIII,IIOOI00000OO00O10l1lOIIIOl1lIOIIII=>IIO00110lO0OI1OOI01011ll0II0IOIIII,IO10O0OI111O0III0OI0Ol0I0llOOIIIII=>II001O10OO10OI0l00lOI0OlOI0IOIIIII,IOOllO1OO0IlII00llll11I1IIO1IIIIII=>
IOlOI0l01llI0OI011lO0010II101IIIII);END GENERATE;S_AXIS_A_TREADY<='1'WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_RATE>1 AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_LATENCY=0)ELSE IOI0l1l111IIIOOO01I0lOO1l1Il0IIIII WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_CE_THROTTLE OR IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_THROTTLE_SCHEME=CI_RFD_THROTTLE OR IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_GEN_THROTTLE OR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=
CI_AND_TVALID_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1))ELSE 'X';S_AXIS_B_TREADY<='1'WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B=1 AND(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1 AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_LATENCY=0))ELSE IO0lI1lO1000O00IO0l00Ol1lOIl1IIIII WHEN(
IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_B=1 AND(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_CE_THROTTLE OR IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE OR
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_GEN_THROTTLE OR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1)))
ELSE 'X';S_AXIS_OPERATION_TREADY<='1'WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION=1 AND(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE AND
 IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1 AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_LATENCY=0))ELSE IOOl010OO0lO0111O00l0Il1I1O1OIIIII WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_OPERATION=1 AND(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII
.C_THROTTLE_SCHEME=CI_CE_THROTTLE OR IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_RFD_THROTTLE OR IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_GEN_THROTTLE
 OR(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_THROTTLE_SCHEME=CI_AND_TVALID_THROTTLE AND IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_RATE>1)))ELSE 'X';M_AXIS_RESULT_TVALID<=
IIO00110IlIOl01O1I0O10100O111IIIII;M_AXIS_RESULT_TDATA<=IIO00110lO0OI1OOI01011ll0II0IOIIII;M_AXIS_RESULT_TUSER<=II001O10OO10OI0l00lOI0OlOI0IOIIIII WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.
C_HAS_RESULT_TUSER=1)ELSE(OTHERS=>'X');M_AXIS_RESULT_TLAST<=IOlOI0l01llI0OI011lO0010II101IIIII WHEN(IOIl10IlOIlOO1lI1lII1llOIIlIOIIIII.C_HAS_RESULT_TLAST=1)ELSE 'X';END
;
