-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /   Vendor: Xilinx
-- \   \   \/    Version: 4.0
--  \   \        Filename: $RCSfile: dds_compiler_v5_0.vhd,v $
--  /   /        Date Last Modified: $Date: 2010/09/08 11:21:20 $
-- /___/   /\    Date Created: 2006
-- \   \  /  \
--  \___\/\___\
--
-- Device  : All
-- Library : dds_compiler_v5_0
-- Purpose : Entity-architecture for XST level core interface
-------------------------------------------------------------------------------
--  (c) Copyright 2006-2010 Xilinx, Inc. All rights reserved.
--
--  This file contains confidential and proprietary information
--  of Xilinx, Inc. and is protected under U.S. and
--  international copyright and other intellectual property
--  laws.
--
--  DISCLAIMER
--  This disclaimer is not a license and does not grant any
--  rights to the materials distributed herewith. Except as
--  otherwise provided in a valid license issued to you by
--  Xilinx, and to the maximum extent permitted by applicable
--  law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
--  WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
--  AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
--  BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
--  INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
--  (2) Xilinx shall not be liable (whether in contract or tort,
--  including negligence, or under any other theory of
--  liability) for any loss or damage of any kind or nature
--  related to, arising under or in connection with these
--  materials, including for any direct, or any indirect,
--  special, incidental, or consequential loss or damage
--  (including loss of data, profits, goodwill, or any type of
--  loss or damage suffered as a result of any action brought
--  by a third party) even if such damage or loss was
--  reasonably foreseeable or Xilinx had been advised of the
--  possibility of the same.
--
--  CRITICAL APPLICATIONS
--  Xilinx products are not designed or intended to be fail-
--  safe, or for use in any application requiring fail-safe
--  performance, such as life-support or safety devices or
--  systems, Class III medical devices, nuclear facilities,
--  applications related to the deployment of airbags, or any
--  other applications that could lead to death, personal
--  injury, or severe property or environmental damage
--  (individually and collectively, "Critical
--  Applications"). Customer assumes the sole risk and
--  liability of any use of Xilinx products in Critical
--  Applications, subject only to applicable laws and
--  regulations governing limitations on product liability.
--
--  THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
--  PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Synthesizable model, AXI-S wrapper
--
-- Adds FIFO logic for AXI interface, instantiates original core as-is with
-- port remapping
--
-- ### WARNING!!!  DO NOT EDIT THIS FILE BY HAND!  USE cp_to_sim.sh IN hdl/ INSTEAD! ###
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library xilinxcorelib;
use xilinxcorelib.pkg_dds_compiler_v5_0.all;
use xilinxcorelib.dds_compiler_v5_0_sim_comps.all;

library xilinxcorelib;
use xilinxcorelib.bip_utils_pkg_v2_0.all;
use xilinxcorelib.xcc_utils_v2_0.all;

library xilinxcorelib;
use xilinxcorelib.xbip_pipe_v2_0_xst_comp.all;

library xilinxcorelib;
use xilinxcorelib.axi_utils_pkg_v1_0.all;
use xilinxcorelib.axi_utils_v1_0_comps.all;

--core_if on entity dds_compiler_v5_0
entity dds_compiler_v5_0 is
  generic (
    C_XDEVICEFAMILY                 :     string                                              := "virtex6";
    C_ACCUMULATOR_WIDTH             :     integer                                             := 28;  -- width of accum and associated paths. Factor in Frequency resolution
    C_CHANNELS                      :     integer                                             := 1;  -- number of time-multiplexed channels output
    C_HAS_CHANNEL_INDEX             :     integer                                             := 0;  -- enables CHANNEL output port
    C_HAS_PHASE_OUT                 :     integer                                             := 0;  -- phase_out pin visible
    C_HAS_PHASEGEN                  :     integer                                             := 1;  -- generate the phase accumulator
    C_HAS_SINCOS                    :     integer                                             := 1;  -- generate the sin/cos block
    C_LATENCY                       :     integer                                             := -1;  -- Selects overall latency, -1 means 'fully pipelined for max performance'
    C_MEM_TYPE                      :     integer                                             := 1;  -- 0= Auto, 1 = Block ROM, 2 = DIST_ROM
    C_NEGATIVE_COSINE               :     integer                                             := 0;  -- 0 = normal cosine, 1 = negated COSINE output port
    C_NEGATIVE_SINE                 :     integer                                             := 0;  -- 0 = normal sine, 1 = negated SINE output port
    C_NOISE_SHAPING                 :     integer                                             := 0;  -- 0 = none, 1 = Dither, 2 = Error Feed Forward (Taylor)
    C_OUTPUTS_REQUIRED              :     integer                                             := 2;  -- 0 = SIN, 1 = COS, 2 = Both;
    C_OUTPUT_WIDTH                  :     integer                                             := 6;  -- sets width of output port (factor in SFDR)
    C_PHASE_ANGLE_WIDTH             :     integer                                             := 6;  -- width of phase fed to RAM (factor in RAM resource used)
    C_PHASE_INCREMENT               :     integer                                             := 2;  -- 1 = register, 2 = constant, 3 = streaming (input port);
    C_PHASE_INCREMENT_VALUE         :     string                                              := "0";  -- string of values for PINC, one for each channel.
    C_PHASE_OFFSET                  :     integer                                             := 0;  -- 0 = none, 1 = reg, 2 = const, 3 = stream (input port);
    C_PHASE_OFFSET_VALUE            :     string                                              := "0";  -- string of values for POFF, one for each channel
    C_OPTIMISE_GOAL                 :     integer                                             := 0;  -- 0 = area, 1 = speed
    C_USE_DSP48                     :     integer                                             := 0;  -- 0 = minimal 1 = max. Determines DSP48 use in phase accumulation.
    C_POR_MODE                      :     integer                                             := 0;  -- Power-on-reset behaviour (for behavioral model)
    C_AMPLITUDE                     :     integer                                             := 0;  -- 0 = full scale (+/- 2^N-2), 1 = unit circle (+/- 2^(N-1))
    -------------------------------------------------------------------------
    -- AXI-S interface generics
    -------------------------------------------------------------------------
    -- General
    C_HAS_ACLKEN                    :     integer                                             := 0;  -- enables active-high clock enable
    C_HAS_ARESETN                   :     integer                                             := 0;  -- enables active-low synchronous reset
    C_HAS_TLAST                     :     integer                                             := 0;  -- enables TLAST signals on relevant channels
    C_HAS_TREADY                    :     integer                                             := 1;  -- enables TREADY signals on relevant channels
    -- S_PHASE
    C_HAS_S_PHASE                   :     integer                                             := 1;  -- enables phase input channel
    C_S_PHASE_TDATA_WIDTH           :     integer                                             := 8;  -- TDATA width (byte-sized)
    C_S_PHASE_HAS_TUSER             :     integer                                             := 0;  -- enables phase channel TUSER, selects TUSER content
    C_S_PHASE_TUSER_WIDTH           :     integer                                             := 1;  -- TUSER width
    -- S_CONFIG
    C_HAS_S_CONFIG                  :     integer                                             := 0;  -- enables config input channel
    C_S_CONFIG_SYNC_MODE            :     integer                                             := 0;  -- specifies how config is synchronized to phase channel
    C_S_CONFIG_TDATA_WIDTH          :     integer                                             := 0;  -- TDATA width (byte-sized)
    -- M_DATA
    C_HAS_M_DATA                    :     integer                                             := 1;  -- enables data output channel
    C_M_DATA_TDATA_WIDTH            :     integer                                             := 32;  -- TDATA width (byte-sized)
    C_M_DATA_HAS_TUSER              :     integer                                             := 0;  -- enables data channel TUSER, selects TUSER content
    C_M_DATA_TUSER_WIDTH            :     integer                                             := 1;  -- TUSER width
    -- M_PHASE
    C_HAS_M_PHASE                   :     integer                                             := 0;  -- enables phase output channel
    C_M_PHASE_TDATA_WIDTH           :     integer                                             := 0;  -- TDATA width (byte-sized)
    C_M_PHASE_HAS_TUSER             :     integer                                             := 0;  -- enables phase channel TUSER, selects TUSER content
    C_M_PHASE_TUSER_WIDTH           :     integer                                             := 1;  -- TUSER width
    ---------------------------------------------------------------------------
    -- Debug/validation enablement
    ---------------------------------------------------------------------------
    C_DEBUG_INTERFACE               :     integer                                             := 0;
    C_CHAN_WIDTH                    :     integer                                             := 1
    );
  port (
    -- Common ports
    aclk                            : in  std_logic                                           := '0';
    aclken                          : in  std_logic                                           := '1';
    aresetn                         : in  std_logic                                           := '1';
    -- S_PHASE
    s_axis_phase_tvalid             : in  std_logic                                           := '0';
    s_axis_phase_tready             : out std_logic                                           := '0';
    s_axis_phase_tdata              : in  std_logic_vector(C_S_PHASE_TDATA_WIDTH-1 downto 0)  := (others => '0');
    s_axis_phase_tlast              : in  std_logic                                           := '0';
    s_axis_phase_tuser              : in  std_logic_vector(C_S_PHASE_TUSER_WIDTH-1 downto 0)  := (others => '0');
    -- S_CONFIG
    s_axis_config_tvalid            : in  std_logic                                           := '0';
    s_axis_config_tready            : out std_logic                                           := '0';
    s_axis_config_tdata             : in  std_logic_vector(C_S_CONFIG_TDATA_WIDTH-1 downto 0) := (others => '0');
    s_axis_config_tlast             : in  std_logic                                           := '0';
    -- M_DATA
    m_axis_data_tvalid              : out std_logic                                           := '0';
    m_axis_data_tready              : in  std_logic                                           := '0';
    m_axis_data_tdata               : out std_logic_vector(C_M_DATA_TDATA_WIDTH-1 downto 0)   := (others => '0');
    m_axis_data_tlast               : out std_logic                                           := '0';
    m_axis_data_tuser               : out std_logic_vector(C_M_DATA_TUSER_WIDTH-1 downto 0)   := (others => '0');
    -- M_PHASE
    m_axis_phase_tvalid             : out std_logic                                           := '0';
    m_axis_phase_tready             : in  std_logic                                           := '0';
    m_axis_phase_tdata              : out std_logic_vector(C_M_PHASE_TDATA_WIDTH-1 downto 0)  := (others => '0');
    m_axis_phase_tlast              : out std_logic                                           := '0';
    m_axis_phase_tuser              : out std_logic_vector(C_M_PHASE_TUSER_WIDTH-1 downto 0)  := (others => '0');
    -- Event Interface
    event_s_phase_tlast_missing     : out std_logic                                           := '0';
    event_s_phase_tlast_unexpected  : out std_logic                                           := '0';
    event_s_phase_chanid_incorrect  : out std_logic                                           := '0';
    event_s_config_tlast_missing    : out std_logic                                           := '0';
    event_s_config_tlast_unexpected : out std_logic                                           := '0';
    -- Debug ports
    debug_axi_pinc_in               : out std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)    := (others => '0');
    debug_axi_poff_in               : out std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)    := (others => '0');
    debug_axi_chan_in               : out std_logic_vector(C_CHAN_WIDTH-1 downto 0)           := (others => '0');
    debug_core_nd                   : out std_logic                                           := '0';
    debug_phase                     : out std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)    := (others => '0');
    debug_phase_nd                  : out std_logic                                           := '0'
    );
--core_if off
end dds_compiler_v5_0;

architecture behavioral of dds_compiler_v5_0 is

  constant singlechannel : boolean := (C_CHANNELS = 1);
  constant multichannel  : boolean := (C_CHANNELS > 1);
  constant lastchannel   : integer := C_CHANNELS-1;

  constant ci_check_generics : integer := check_generics(
    P_XDEVICEFAMILY         => C_XDEVICEFAMILY,
    P_ACCUMULATOR_WIDTH     => C_ACCUMULATOR_WIDTH,
    P_CHANNELS              => C_CHANNELS,
    P_HAS_CHANNEL_INDEX     => C_HAS_CHANNEL_INDEX,
    P_HAS_PHASE_OUT         => C_HAS_PHASE_OUT,
    P_HAS_PHASEGEN          => C_HAS_PHASEGEN,
    P_HAS_SINCOS            => C_HAS_SINCOS,
    P_LATENCY               => C_LATENCY,
    P_MEM_TYPE              => C_MEM_TYPE,
    P_NEGATIVE_COSINE       => C_NEGATIVE_COSINE,
    P_NEGATIVE_SINE         => C_NEGATIVE_SINE,
    P_NOISE_SHAPING         => C_NOISE_SHAPING,
    P_OUTPUTS_REQUIRED      => C_OUTPUTS_REQUIRED,
    P_OUTPUT_WIDTH          => C_OUTPUT_WIDTH,
    P_PHASE_ANGLE_WIDTH     => C_PHASE_ANGLE_WIDTH,
    P_PHASE_INCREMENT       => C_PHASE_INCREMENT,
    P_PHASE_INCREMENT_VALUE => C_PHASE_INCREMENT_VALUE,
    P_PHASE_OFFSET          => C_PHASE_OFFSET,
    P_PHASE_OFFSET_VALUE    => C_PHASE_OFFSET_VALUE,
    P_OPTIMISE_GOAL         => C_OPTIMISE_GOAL,
    P_USE_DSP48             => C_USE_DSP48,
    P_POR_MODE              => C_POR_MODE,
    P_AMPLITUDE             => C_AMPLITUDE,
    -- General
    P_HAS_ACLKEN            => C_HAS_ACLKEN,
    P_HAS_ARESETN           => C_HAS_ARESETN,
    P_HAS_TLAST             => C_HAS_TLAST,
    P_HAS_TREADY            => C_HAS_TREADY,
    -- S_PHASE
    P_HAS_S_PHASE           => C_HAS_S_PHASE,
    P_S_PHASE_TDATA_WIDTH   => C_S_PHASE_TDATA_WIDTH,
    P_S_PHASE_HAS_TUSER     => C_S_PHASE_HAS_TUSER,
    P_S_PHASE_TUSER_WIDTH   => C_S_PHASE_TUSER_WIDTH,
    -- S_CONFIG
    P_HAS_S_CONFIG          => C_HAS_S_CONFIG,
    P_S_CONFIG_SYNC_MODE    => C_S_CONFIG_SYNC_MODE,
    P_S_CONFIG_TDATA_WIDTH  => C_S_CONFIG_TDATA_WIDTH,
    -- M_DATA
    P_HAS_M_DATA            => C_HAS_M_DATA,
    P_M_DATA_TDATA_WIDTH    => C_M_DATA_TDATA_WIDTH,
    P_M_DATA_HAS_TUSER      => C_M_DATA_HAS_TUSER,
    P_M_DATA_TUSER_WIDTH    => C_M_DATA_TUSER_WIDTH,
    -- M_PHASE
    P_HAS_M_PHASE           => C_HAS_M_PHASE,
    P_M_PHASE_TDATA_WIDTH   => C_M_PHASE_TDATA_WIDTH,
    P_M_PHASE_HAS_TUSER     => C_M_PHASE_HAS_TUSER,
    P_M_PHASE_TUSER_WIDTH   => C_M_PHASE_TUSER_WIDTH
    );

  constant ci_axi_latency_overhead   : integer := fn_get_axi_latency_overhead(
    p_has_tready      => C_HAS_TREADY,
    p_phase_increment => C_PHASE_INCREMENT,
    p_phase_offset    => C_PHASE_OFFSET
    );
  signal   diag_axi_latency_overhead : integer := ci_axi_latency_overhead;

  constant ci_core_latency   : integer := fn_get_core_latency(
    p_axi_overhead => ci_axi_latency_overhead,
    p_latency      => C_LATENCY
    );
  signal   diag_core_latency : integer := ci_core_latency;

  signal sclr_i   : std_logic := '0';
  signal aclken_i : std_logic := '1';

  signal ce_i, ce_i_delayed, ce_core : std_logic := '0';

  -- Delay between asking for a read, and getting the data back
  constant srl_fifo_turnaround_latency : integer := 1;

  -----------------------------------------------------------------------------
  -- Important note. Internal, legacy core is configured to take inputs from
  -- AXI or not. When it does, the internal core is set to streaming and all
  -- inputs generated from AXI interface. When not (source-only), the core can
  -- produce its own channel out, RDY, etc.
  -----------------------------------------------------------------------------
  constant ci_int_core_mode : t_int_core_mode := fn_resolve_int_core_mode(
    p_channels        => C_CHANNELS,
    p_has_phase_gen   => C_HAS_PHASEGEN,
    p_phase_increment => C_PHASE_INCREMENT,
    p_phase_offset    => C_PHASE_OFFSET
    );

  signal diag_int_core_mode : t_int_core_mode := ci_int_core_mode;

  constant dds_latencies : t_latency_allocation_return := fn_dds_compiler_v5_0_latency(
    p_xdevicefamily     => C_XDEVICEFAMILY,
    p_has_phasegen      => C_HAS_PHASEGEN,
    p_has_sincos        => C_HAS_SINCOS,
    p_latency           => ci_core_latency,  -- NOTE: not C_LATENCY!
    p_mem_type          => C_MEM_TYPE,
    p_accumulator_width => C_ACCUMULATOR_WIDTH,
    p_noise_shaping     => C_NOISE_SHAPING,
    p_phase_angle_width => C_PHASE_ANGLE_WIDTH,
    p_phase_increment   => ci_int_core_mode.phase_inc,
    p_phase_offset      => ci_int_core_mode.phase_offset,
    p_optimise_goal     => C_OPTIMISE_GOAL,
    p_use_dsp48         => C_USE_DSP48,
    p_channels          => C_CHANNELS,
    p_output_width      => C_OUTPUT_WIDTH
    );

  constant dds_pipeline_latency  : integer := dds_latencies.used;
  constant dds_sincos_latency    : integer := dds_latencies.sc_lat;
  constant dds_phase_gen_latency : integer := dds_latencies.pg_lat;
  constant dds_lump1_latency     : integer := dds_latencies.lump_lat_1;
  constant dds_lump2_latency     : integer := dds_latencies.lump_lat_2;

  constant ci_dither_delay : t_dither_delays := fn_dither_delay(
    p_pipe            => dds_latencies.pipe,
    p_use_dsp48       => fn_use_dsp48(C_USE_DSP48, C_XDEVICEFAMILY),
    p_xdevicefamily   => C_XDEVICEFAMILY,
    p_channels        => C_CHANNELS,
    p_phase_increment => C_PHASE_INCREMENT,
    p_phase_offset    => C_PHASE_OFFSET
    );

  constant dds_dither_delay : integer := ci_dither_delay.datapath;


-- For latency debug
-- function report_lat
-- return integer is
-- begin
-- report "dds_pipeline_latency " & integer'image(dds_pipeline_latency) severity note;
-- report "dds_sincos_latency " & integer'image(dds_sincos_latency) severity note;
-- report "dds_phase_gen_latency " & integer'image(dds_phase_gen_latency) severity note;
-- report "dds_lump1 latency " & integer'image(dds_latencies.lump_lat_1) severity note;
-- report "dds_lump2_latency " & integer'image(dds_latencies.lump_lat_2) severity note;
-- report "dither datapath lat " & integer'image(dds_dither_delay) severity note;
-- return 0;
-- end function report_lat;
-- constant get_lat : integer := report_lat;

  signal nd_i, rdy_stream_i : std_logic := '0';

  constant ci_chan_width : integer := sel_lines_reqd(C_CHANNELS);

  constant ci_phase_inc_inits     : t_ram_type                                       := fn_init_ram(C_PHASE_INCREMENT_VALUE, C_CHANNELS, ci_chan_width, C_ACCUMULATOR_WIDTH);
  constant ci_phase_adj_inits     : t_ram_type                                       := fn_init_ram(C_PHASE_OFFSET_VALUE, C_CHANNELS, ci_chan_width, C_ACCUMULATOR_WIDTH);
  constant ci_phase_inc_acc_inits : t_ram_type                                       := fn_init_ram(C_PHASE_INCREMENT_VALUE, C_CHANNELS, ci_chan_width, C_ACCUMULATOR_WIDTH);
  constant ci_phase_adj_acc_inits : t_ram_type                                       := fn_init_ram(C_PHASE_OFFSET_VALUE, C_CHANNELS, ci_chan_width, C_ACCUMULATOR_WIDTH);
  constant ci_phase_inc           : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := ci_phase_inc_acc_inits(0)(C_ACCUMULATOR_WIDTH-1 downto 0);
  constant ci_phase_adj           : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := ci_phase_adj_acc_inits(0)(C_ACCUMULATOR_WIDTH-1 downto 0);
  signal   diag_phase_inc_inits   : t_ram_type                                       := ci_phase_inc_inits;
  signal   diag_phase_adj_inits   : t_ram_type                                       := ci_phase_adj_inits;

  -----------------------------------------------------------------------------
  -- DDS internal core signals
  -----------------------------------------------------------------------------
  signal dds_pinc_in : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
  signal dds_poff_in : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
  signal dds_rdy     : std_logic                                        := '0';

  --When the old core is configured as source, use it's output channel
  --When the old core is configured as a streamer, use the AXI input channel count.
  --Whichever you use, call it dds_channel.
  signal dds_channel         : std_logic_vector(ci_chan_width-1 downto 0) := (others => '0');
  signal legacy_core_channel : std_logic_vector(ci_chan_width-1 downto 0) := (others => '0');
  signal stream_channel      : std_logic_vector(ci_chan_width-1 downto 0) := (others => '0');

  signal dds_cosine    : std_logic_vector(C_OUTPUT_WIDTH-1 downto 0)      := (others => '0');
  signal dds_sine      : std_logic_vector(C_OUTPUT_WIDTH-1 downto 0)      := (others => '0');
  signal dds_phase_out : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');

  signal   dds_addr                     : std_logic_vector(sel_lines_reqd(C_CHANNELS)-1 downto 0) := (others => '0');
  constant dds_reg_select_dummy         : std_logic                                               := '0';
  signal   dds_we                       : std_logic                                               := '0';
  constant dds_data_dummy               : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)        := (others => '0');
  signal   dds_pinc_data, dds_poff_data : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)        := (others => '0');
  signal   dds_debug_phase              : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0)        := (others => '0');

  -----------------------------------------------------------------------------
  -- Signals for input FIFOs
  -----------------------------------------------------------------------------
  constant s_phase_fifo_width                                                                                         : integer                                         := calc_s_phase_fifo_width(C_HAS_PHASEGEN, C_ACCUMULATOR_WIDTH, C_PHASE_INCREMENT, C_PHASE_OFFSET, C_S_PHASE_HAS_TUSER, C_S_PHASE_TUSER_WIDTH, C_HAS_TLAST, C_CHANNELS);
  signal   s_phase_fifo_din, s_phase_fifo_dout                                                                        : std_logic_vector(s_phase_fifo_width-1 downto 0) := (others => '0');
  signal   s_phase_fifo_rd_enable, s_phase_fifo_rd_avail, s_phase_fifo_rd_valid, s_phase_fifo_not_empty               : std_logic                                       := '0';
  signal   s_phase_tlast                                                                                              : std_logic                                       := '0';
  -- for debug
  signal   s_phase_fifo_full, s_phase_fifo_empty, s_phase_fifo_aempty, s_phase_fifo_not_full, s_phase_fifo_not_aempty : std_logic                                       := '0';
  signal   s_phase_fifo_add                                                                                           : signed(4 downto 0)                              := (others => '0');

  signal chanid_in         : std_logic_vector(sel_lines_reqd(C_CHANNELS)-1 downto 0);
  signal user_in, user_out : std_logic_vector(calc_user_in_width(C_CHANNELS, C_S_PHASE_HAS_TUSER, C_S_PHASE_TUSER_WIDTH, C_HAS_TLAST)-1 downto 0);

  signal s_axis_config_tready_pre : std_logic := '0';
  signal s_axis_config_tready_i   : std_logic := '0';
  -----------------------------------------------------------------------------
  -- Signals for output FIFOs
  -----------------------------------------------------------------------------

  constant m_data_fifo_width                                         : integer                                        := calc_m_data_fifo_width(C_OUTPUT_WIDTH, C_OUTPUTS_REQUIRED, C_M_DATA_HAS_TUSER, C_M_DATA_TUSER_WIDTH, C_HAS_TLAST);
  constant m_data_fifo_depth                                         : integer                                        := 16;
  signal   m_data_fifo_din, m_data_fifo_dout                         : std_logic_vector(m_data_fifo_width-1 downto 0) := (others => '0');
  signal   m_data_fifo_wr_enable                                     : std_logic                                      := '0';
  signal   m_data_fifo_not_afull                                     : std_logic                                      := '1';
  -- for debug
  signal   m_data_fifo_full, m_data_fifo_afull, m_data_fifo_not_full : std_logic                                      := '0';

  constant m_phase_fifo_width                                           : integer                                         := calc_m_phase_fifo_width(C_ACCUMULATOR_WIDTH, C_M_PHASE_HAS_TUSER, C_M_PHASE_TUSER_WIDTH, C_HAS_TLAST);
  constant m_phase_fifo_depth                                           : integer                                         := 16;
  signal   m_phase_fifo_din, m_phase_fifo_dout                          : std_logic_vector(m_phase_fifo_width-1 downto 0) := (others => '0');
  signal   m_phase_fifo_wr_enable                                       : std_logic                                       := '0';
  signal   m_phase_fifo_not_afull                                       : std_logic                                       := '1';
  -- for debug
  signal   m_phase_fifo_full, m_phase_fifo_afull, m_phase_fifo_not_full : std_logic                                       := '0';

  signal pull_data : std_logic := '0';

  constant dds_cfg : R_DDS_CFG := (
    outputs_required     => C_OUTPUTS_REQUIRED,
    has_phase_out        => C_HAS_PHASE_OUT,
    output_width         => C_OUTPUT_WIDTH,
    channels             => C_CHANNELS,
    has_phasegen         => C_HAS_PHASEGEN,
    has_sincos           => C_HAS_SINCOS,
    phase_increment      => C_PHASE_INCREMENT,
    phase_offset         => C_PHASE_OFFSET,
    accumulator_width    => C_ACCUMULATOR_WIDTH,
    has_tlast            => C_HAS_TLAST,
    has_s_config         => C_HAS_S_CONFIG,
    has_s_phase          => C_HAS_S_PHASE,
    has_m_data           => C_HAS_M_DATA,
    has_m_phase          => C_HAS_M_PHASE,
    s_config_tdata_width => C_S_CONFIG_TDATA_WIDTH,
    s_phase_tdata_width  => C_S_PHASE_TDATA_WIDTH,
    s_phase_has_tuser    => C_S_PHASE_HAS_TUSER,
    s_phase_tuser_width  => C_S_PHASE_TUSER_WIDTH,
    m_data_tdata_width   => C_M_DATA_TDATA_WIDTH,
    m_data_has_tuser     => C_M_DATA_HAS_TUSER,
    m_data_tuser_width   => C_M_DATA_TUSER_WIDTH,
    m_phase_tdata_width  => C_M_PHASE_TDATA_WIDTH,
    m_phase_has_tuser    => C_M_PHASE_HAS_TUSER,
    m_phase_tuser_width  => C_M_PHASE_TUSER_WIDTH
    );

  signal addr_counter     : unsigned(sel_lines_reqd(C_CHANNELS)-1 downto 0) := (others => '0');
  signal addr_counter_max : std_logic                                       := '0';

  signal tlast_out : std_logic := '0';

  --diagnostic loom signals - datum for validation. These signals demark the
  --end of the input circuitry and the start of the legacy DDS.
  signal axi_pinc_in  : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
  signal axi_poff_in  : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
  signal axi_phase_in : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
  signal axi_chan_in  : std_logic_vector(ci_chan_width-1 downto 0)       := (others => '0');
  signal axi_tlast_in : std_logic                                        := '0';

  signal   master_count     : unsigned(ci_chan_width-1 downto 0) := (others => '0');  --master channel counter
  constant master_count_inc : unsigned(ci_chan_width-1 downto 0) := to_unsigned(1, ci_chan_width);  --long way round to say "+1"

begin

  -----------------------------------------------------------------------------
  -- Set up common signals
  -----------------------------------------------------------------------------

  has_aclken : if C_HAS_ACLKEN = 1 generate
    aclken_i <= aclken;
  end generate has_aclken;

  has_aresetn             : if C_HAS_ARESETN = 1 generate
    signal reset_history  : std_logic_vector(2 downto 0) := (others => '0');
  begin
    sclr_i_reg            : process (aclk) is
    begin
      if rising_edge(aclk) then
        sclr_i        <= not aresetn;
      end if;
    end process sclr_i_reg;
    -- synthesis translate_off
    check_reset           : process (aclk) is
    begin
      if rising_edge(aclk) then
        reset_history <= reset_history(1 downto 0) & ARESETN;
        assert not(reset_history = "010" or reset_history = "101")
          report "WARNING : aresetn must be asserted or deasserted for a minimum of 2 cycles"
          severity warning;
      end if;
    end process check_reset;
    -- synthesis translate_on
  end generate has_aresetn;

  -- Enable for DDS sub-module so pipeline is stalled when
  ce_i <= aclken_i and pull_data;



  --This is the nd-rdy pipeline.
  i_has_nd_rdy_pipe      : if ci_int_core_mode.int_core = ci_int_core_mode_streaming generate
    valid_phase_read_del : xbip_pipe_v2_0_xst
      generic map(
        C_LATENCY  => dds_pipeline_latency,
        C_HAS_CE   => 1,
        C_HAS_SCLR => 1,
        C_WIDTH    => 1
        )
      port map(
        CLK        => aclk,
        CE         => ce_core,
        SCLR       => sclr_i,
        D(0)       => nd_i,
        Q(0)       => rdy_stream_i
        );
    channel_pipe         : xbip_pipe_v2_0_xst
      generic map(
        C_LATENCY  => dds_pipeline_latency,
        C_HAS_CE   => 1,
        C_HAS_SCLR => 1,
        C_WIDTH    => ci_chan_width
        )
      port map(
        CLK        => aclk,
        CE         => ce_core,
        SCLR       => sclr_i,
        D          => axi_chan_in,
        Q          => stream_channel
        );
  end generate i_has_nd_rdy_pipe;

  nd_i    <= ce_core;

  i_has_no_phase : if C_HAS_S_PHASE = 0 generate
    ce_core <= ce_i;
  end generate i_has_no_phase;
  -----------------------------------------------------------------------------
  -- CE selection
  -----------------------------------------------------------------------------
  i_ce_s_phase : if C_HAS_S_PHASE = 1 generate
    i_has_tready : if C_HAS_TREADY = 1 generate
      ce_core <= ce_i_delayed and s_phase_fifo_rd_valid;
    end generate i_has_tready;
    i_has_no_tready : if C_HAS_TREADY = 0 generate
      -- We don't do bubble insertion.  We effectively push data through the
      -- core when there's no ready
      ce_core <= ce_i and (s_axis_phase_tvalid and aclken_i);
    end generate i_has_no_tready;
  end generate i_ce_s_phase;

  has_s_phase : if C_HAS_S_PHASE = 1 generate

    s_phase_fifo_din(s_phase_fifo_width-1 downto 0) <= build_s_phase_fifo_din (
      dds_cfg,
      s_phase_fifo_width,
      s_axis_phase_tdata,
      s_axis_phase_tuser,
      s_axis_phase_tlast
      );

    i_with_tready  : if C_HAS_TREADY = 1 generate
      s_phase_fifo : glb_ifx_slave_v1_0
        generic map(
          WIDTH          => s_phase_fifo_width,
          DEPTH          => 16,
          HAS_UVPROT     => true,
          HAS_IFX        => false,
          AEMPTY_THRESH0 => 0,
          AEMPTY_THRESH1 => 0
          )
        port map(
          aclk           => aclk,
          aclken         => aclken_i,
          areset         => sclr_i,     -- REVISIT: not need to reset instantly?
          ifx_valid      => s_axis_phase_tvalid,
          ifx_ready      => s_axis_phase_tready,
          ifx_data       => s_phase_fifo_din,
          -- read interface
          rd_enable      => s_phase_fifo_rd_enable,
          rd_avail       => s_phase_fifo_rd_avail,
          rd_valid       => s_phase_fifo_rd_valid,
          rd_data        => s_phase_fifo_dout,
          -- status
          full           => s_phase_fifo_full,
          empty          => s_phase_fifo_empty,
          aempty         => s_phase_fifo_aempty,
          not_full       => s_phase_fifo_not_full,
          not_empty      => s_phase_fifo_not_empty,
          not_aempty     => s_phase_fifo_not_aempty,
          add            => s_phase_fifo_add
          );

      s_phase_fifo_rd_enable <= ce_i and s_phase_fifo_rd_avail;

    end generate i_with_tready;

    i_has_no_tready               : if C_HAS_TREADY = 0 generate
      signal reg_s_phase_fifo_din : std_logic_vector(s_phase_fifo_width-1 downto 0) := (others => '0');
    begin
      s_phase_fifo_dout          <= s_phase_fifo_din when s_axis_phase_tvalid = '1' else reg_s_phase_fifo_din;
      i_s_phase_halfaxi_reg       : process(aclk)
      begin
        if rising_edge(aclk) then
          if sclr_i = '1' then
            reg_s_phase_fifo_din <= (others                                                    => '0');
          elsif aclken_i = '1' then
            reg_s_phase_fifo_din <= s_phase_fifo_dout;
          end if;
        end if;
      end process i_s_phase_halfaxi_reg;
    end generate i_has_no_tready;

    -- only need to delay internal CE to core when FIFO is present
    ce_i_delay : xbip_pipe_v2_0_xst
      generic map(
        C_LATENCY  => srl_fifo_turnaround_latency,
        C_HAS_CE   => C_HAS_ACLKEN,
        C_HAS_SCLR => 1,
        C_WIDTH    => 1
        )
      port map(
        CLK        => aclk,
        CE         => '1',
        SCLR       => sclr_i,
        D(0)       => ce_i,
        Q(0)       => ce_i_delayed
        );

    decompose_s_phase_fifo_dout (
      dds_cfg            => dds_cfg,
      s_phase_fifo_width => s_phase_fifo_width,
      s_phase_fifo_dout  => s_phase_fifo_dout,
      pinc               => dds_pinc_in,
      poff               => dds_poff_in,
      phase_in           => axi_phase_in,
      chanid             => chanid_in,
      user               => user_in,
      tlast              => s_phase_tlast);


    -- Build TUSER delay
    has_input_tuser : if C_S_PHASE_HAS_TUSER = ci_tuser_user_field or C_S_PHASE_HAS_TUSER = ci_tuser_user_field_and_chanid generate
      -- No reset required as outputs are qualified with TVALID or FIFO write enable
      tuser_delay   : xbip_pipe_v2_0_xst
        generic map(
          C_LATENCY  => dds_pipeline_latency,
          C_HAS_CE   => 1,
          C_HAS_SCLR => 0,
          C_WIDTH    => user_in'length
          )
        port map(
          CLK        => aclk,
          CE         => ce_core,
          SCLR       => '0',
          D          => user_in,
          Q          => user_out
          );
    end generate has_input_tuser;

    -- Event interface
    s_phase_tlast_checks : if C_S_CONFIG_SYNC_MODE = ci_s_config_sync_mode_vector generate
      tlast_compare      : process (aclk) is
      begin
        if rising_edge(aclk) then
          if ce_core = '1' then
            if master_count = to_unsigned(lastchannel, master_count'length) then
              -- Reached last channel, but didn't see a TLAST
              event_s_phase_tlast_missing    <= not(s_phase_tlast);
              event_s_phase_tlast_unexpected <= '0';
            else
              event_s_phase_tlast_missing    <= '0';
              -- Didn't reach last channel yet, but got a TLAST for some reason
              event_s_phase_tlast_unexpected <= s_phase_tlast;
            end if;
          end if;
        end if;
      end process tlast_compare;
    end generate s_phase_tlast_checks;

    s_phase_chanid_checks : if C_S_PHASE_HAS_TUSER = ci_tuser_chanid
                              or C_S_PHASE_HAS_TUSER = ci_tuser_user_field_and_chanid generate
      chanid_compare      : process (aclk) is
      begin
        if rising_edge(aclk) then
          if ce_core = '1' then
            if unsigned(chanid_in) /= master_count then
              -- User's channel id didn't match the core's current channel
              event_s_phase_chanid_incorrect <= '1';
            else
              event_s_phase_chanid_incorrect <= '0';
            end if;
          end if;
        end if;
      end process chanid_compare;
    end generate s_phase_chanid_checks;

  end generate has_s_phase;


  -----------------------------------------------------------------------------
  -- Shared master channel count into DDS.
  -----------------------------------------------------------------------------
  master_channel_count : if multichannel generate
    i_master_count     : process(aclk)
    begin
      if rising_edge(aclk) then
        if sclr_i = '1' then
          master_count   <= (others => '0');
        elsif ce_core = '1' then
          if master_count = to_unsigned((lastchannel), master_count'length) then
            master_count <= (others => '0');
          else
            master_count <= master_count + master_count_inc;
          end if;
        end if;
      end if;
    end process i_master_count;
  end generate master_channel_count;



  i_pinc_poff_in                  : if C_HAS_PHASEGEN = 1 generate
    signal   pingpong             : std_logic                                    := '0';
    signal   pingpong_pre         : std_logic                                    := '0';
    signal   config_read_addr     : std_logic_vector(ci_chan_width+1-1 downto 0) := (others => '0');
    signal   config_write_addr    : std_logic_vector(ci_chan_width+1-1 downto 0) := (others => '0');
    signal   config_chan_expected : unsigned(ci_chan_width-1 downto 0)           := (others => '0');  --master channel counter
    constant ci_byte_accum_width  : integer                                      := roundup_to_multiple(C_ACCUMULATOR_WIDTH, 8);
  begin



    s_axis_config_tready         <= s_axis_config_tready_i;
    i_config_multichan       : if multichannel and (C_PHASE_INCREMENT = c_phase_inc_prog or C_PHASE_OFFSET = c_phase_adj_prog) generate
      i_config_chan_expected : process(aclk)
      begin
        if rising_edge(aclk) then
          if sclr_i = '1' then
            config_chan_expected <= (others => '0');
            --else if valid config_write
          elsif s_axis_config_tvalid = '1' and s_axis_config_tready_i = '1' and aclken_i = '1' then

            if config_chan_expected = to_unsigned(lastchannel, config_chan_expected'length) then
              config_chan_expected <= (others => '0');
            else
              config_chan_expected <= config_chan_expected + master_count_inc;
            end if;

            -- Config channel event interface - detect loss of sync when multichannel
--            if C_HAS_TLAST = ci_tlast_vector_framing then. The config channel
--            is ALWAYS vector based.
            if config_chan_expected = to_unsigned(lastchannel, config_chan_expected'length) then
              -- Reached last channel, but didn't see a TLAST
              event_s_config_tlast_missing    <= not(s_axis_config_tlast);
              event_s_config_tlast_unexpected <= '0';
            else
              event_s_config_tlast_missing    <= '0';
              -- Didn't reach last channel yet, but got a TLAST for some reason
              event_s_config_tlast_unexpected <= s_axis_config_tlast;
            end if;
-- end if;                              --not need for if vector based because it's always vector based.

          end if;
        end if;
      end process i_config_chan_expected;
      i_pingpong_reg : xbip_pipe_v2_0_xst
        generic map(
          C_LATENCY  => 1,
          C_HAS_CE   => 1,
          C_HAS_SCLR => 0,
          C_WIDTH    => 1
          )
        port map(
          CLK        => aclk,
          CE         => ce_core,
          SCLR       => '0',            --Note that any valid reconfigurations
          --will survive ARESETN. The power-on init values are lost.
          D(0)       => pingpong_pre,
          Q(0)       => pingpong
          );
      config_write_addr <= not(pingpong) & std_logic_vector(config_chan_expected);
      config_read_addr  <= pingpong & std_logic_vector(master_count);  --REVISIT - needs master channel count.

      --s_axis_config_tready goes low when the input RAM is full goes high on
      --event that toggles pingpong
      i_reconfig_vector_based : if C_S_CONFIG_SYNC_MODE = ci_s_config_sync_mode_vector generate
        s_axis_config_tready_pre <= '1'           when (to_integer(unsigned(config_read_addr(ci_chan_width-1 downto 0))) = lastchannel) and ce_core = '1'                                              else
                                    '0'           when s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel else
                                    s_axis_config_tready_i;
        pingpong_pre             <= not(pingpong) when
                        --trigger moment
                        ((to_integer(unsigned(config_read_addr(ci_chan_width-1 downto 0))) = lastchannel) and ce_core = '1') and
                        --and (been filled
                        (s_axis_config_tready_i = '0' or
                         -- or just filled)
                         (s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel))                            else
                        pingpong;
      end generate i_reconfig_vector_based;
      i_reconfig_packet_based : if C_S_CONFIG_SYNC_MODE = ci_s_config_sync_mode_packet generate
        s_axis_config_tready_pre <= '1'           when (s_phase_tlast = '1') and ce_core = '1'                                                                                                         else
                                    '0'           when s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel else
                                    s_axis_config_tready_i;
        pingpong_pre             <= not(pingpong) when
                        --trigger moment
                        ((s_phase_tlast = '1') and ce_core = '1') and
                        --and (been filled
                        (s_axis_config_tready_i = '0' or
                         -- or just filled)
                         (s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel))                            else
                        pingpong;
      end generate i_reconfig_packet_based;
      i_config_tready_reg     : xbip_pipe_v2_0_xst
        generic map(
          C_LATENCY   => 1,
          C_HAS_CE    => C_HAS_ACLKEN,
          C_HAS_SINIT => 1,
          C_WIDTH     => 1,
          C_SINIT_VAL => "1"
          )
        port map(
          CLK         => aclk,
          CE          => aclken_i,
          SINIT       => sclr_i,
          D(0)        => s_axis_config_tready_pre,
          Q(0)        => s_axis_config_tready_i
          );

      --In this case TLAST means 'last cycle of old configuration', so hold on tight.
      tlast_out_config_triggered_generation : if C_HAS_TLAST = ci_tlast_config_triggered generate
        i_reconfig_vector_based             : if C_S_CONFIG_SYNC_MODE = ci_s_config_sync_mode_vector generate
          axi_tlast_in <= '1' when
                          --trigger moment
                          ((to_integer(unsigned(config_read_addr(ci_chan_width-1 downto 0))) = lastchannel) and ce_core = '1') and
                          --and (been filled
                          (s_axis_config_tready_i = '0' or
                           -- or just filled)
                           (s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel)) else
                          '0';
        end generate i_reconfig_vector_based;
        i_reconfig_packet_based             : if C_S_CONFIG_SYNC_MODE = ci_s_config_sync_mode_packet generate
          axi_tlast_in <= '1' when
                          --trigger moment
                          ((s_phase_tlast = '1') and ce_core = '1') and
                          --and (been filled
                          (s_axis_config_tready_i = '0' or
                           -- or just filled)
                           (s_axis_config_tready_i = '1' and s_axis_config_tvalid = '1' and to_integer(unsigned(config_write_addr(ci_chan_width-1 downto 0))) = lastchannel)) else
                          '0';
        end generate i_reconfig_packet_based;
      end generate tlast_out_config_triggered_generation;

    end generate i_config_multichan;

    i_tready_single_config : if singlechannel and (C_PHASE_INCREMENT = c_phase_inc_prog or C_PHASE_OFFSET = c_phase_adj_prog) generate
      s_axis_config_tready_i <= '1';
    end generate i_tready_single_config;

    -----------------------------------------------------------------------------
    -- Creating fixed, prog and stream input types for PINC
    -- if/generate
    -----------------------------------------------------------------------------
    -- Fixed, single channel.
    i_single_channel_fixed_pinc : if singlechannel and C_PHASE_INCREMENT = c_phase_inc_fixed generate
      axi_pinc_in <= ci_phase_inc;
    end generate i_single_channel_fixed_pinc;

    --Prog, single channel.
    i_single_channel_prog_pinc : if singlechannel and C_PHASE_INCREMENT = c_phase_inc_prog generate
      signal reg_pinc          : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := ci_phase_inc;
      signal config_pinc       : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
    begin
      config_pinc    <= s_axis_config_tdata(C_ACCUMULATOR_WIDTH-1 downto 0);  --this one never moves
      axi_pinc_in    <= config_pinc when s_axis_config_tvalid = '1' else reg_pinc;
      i_pinc_config_reg        : process(aclk)
      begin
        if rising_edge(aclk) then
          if sclr_i = '1' then
            reg_pinc <= ci_phase_inc;
          elsif aclken_i = '1' then
            reg_pinc <= axi_pinc_in;
          end if;
        end if;
      end process i_pinc_config_reg;
    end generate i_single_channel_prog_pinc;

    --Stream, single channel
    i_single_or_mult_channel_stream_pinc : if C_PHASE_INCREMENT = c_phase_inc_streaming generate
      axi_pinc_in <= dds_pinc_in;
    end generate i_single_or_mult_channel_stream_pinc;

    --fixed, Multichannel
    i_mult_channel_fixed_pinc : if multichannel and C_PHASE_INCREMENT = c_phase_inc_fixed generate
      i_inc_ram               : dds_compiler_v5_0_lut_ram
        generic map(
          INIT_VAL     => ci_phase_inc_inits,
          C_CHANNELS   => C_CHANNELS,
          C_DATA_WIDTH => C_ACCUMULATOR_WIDTH,
          C_ADDR_WIDTH => 4,            --unnecessary, but harmless.
          C_DPRA_WIDTH => ci_chan_width,
          C_HAS_MUTE   => 1,            -- contains initial values, so mute always required
          C_HAS_CE     => 1,
          C_LATENCY    => 0
          )
        port map(
          CLK          => aclk,
          --port A
          WE           => '0',
          MUTE         => '0',          --mute_chan, REVISIT G.Old. Needs thought.
          --port B
          CE           => ce_core,
          DPRA         => std_logic_vector(master_count),
          DPO          => axi_pinc_in
          );

    end generate i_mult_channel_fixed_pinc;
    --Prog, Multichannel
    i_mult_channel_prog_pinc : if multichannel and C_PHASE_INCREMENT = c_phase_inc_prog generate
    begin
      i_inc_ram              : dds_compiler_v5_0_lut5_ram
        generic map(
          INIT_VAL     => ci_phase_inc_inits,
          C_CHANNELS   => C_CHANNELS,
          C_DATA_WIDTH => C_ACCUMULATOR_WIDTH,
          C_ADDR_WIDTH => config_write_addr'length,
          C_DPRA_WIDTH => config_read_addr'length,
          C_HAS_MUTE   => 1,            -- contains initial values, so mute always required
          C_HAS_CE     => 1,
          C_LATENCY    => 0             -- allows config to match stream TDM channel
          )
        port map(
          CLK          => aclk,
          --Write side
          WE           => s_axis_config_tvalid,  --REVISIT. and aclken and tready
          --omitted - just let location be overwitten. Last write will be the valid one.
          MUTE         => '0',          --mute_chan,REVISIT - needs thought (as per if gen above)
          A            => config_write_addr,
          DI           => s_axis_config_tdata(C_ACCUMULATOR_WIDTH-1 downto 0),
          --Read side
          CE           => ce_core,
          DPRA         => config_read_addr,  --REVISIT - needs channel addr.
          DPO          => axi_pinc_in
          );

    end generate i_mult_channel_prog_pinc;

    ---------------------------------------------------------------------------
    -- Diag loom addition
    ---------------------------------------------------------------------------
    axi_chan_in   <= std_logic_vector(master_count);  --REVISIT if zero latency master count
                                        --scheme is too slow.
    -----------------------------------------------------------------------------
    -- Creating fixed, prog and stream input types for POFF
    -- if/generate
    -----------------------------------------------------------------------------
    -- Fixed, single channel.
    i_single_channel_fixed_poff : if singlechannel and C_PHASE_OFFSET = c_phase_inc_fixed generate
      axi_poff_in <= ci_phase_adj;
    end generate i_single_channel_fixed_poff;

    --Prog, single channel.
    i_single_channel_prog_poff : if singlechannel and C_PHASE_OFFSET = c_phase_adj_prog generate
      signal pre_reg_poff      : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := ci_phase_adj;
      signal reg_poff          : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := ci_phase_adj;
      signal config_poff       : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
    begin
      --no, really PHASE_INCREMENT
      i_poff_in_upper_tdata    : if C_PHASE_INCREMENT = c_phase_inc_prog generate
        config_poff  <= s_axis_config_tdata(C_ACCUMULATOR_WIDTH + ci_byte_accum_width -1 downto ci_byte_accum_width);
      end generate i_poff_in_upper_tdata;
      --no, really PHASE_INCREMENT
      i_poff_in_lower_tdata    : if C_PHASE_INCREMENT /= c_phase_inc_prog generate  --
        config_poff  <= s_axis_config_tdata(C_ACCUMULATOR_WIDTH-1 downto 0);
      end generate i_poff_in_lower_tdata;
      axi_poff_in    <= config_poff when s_axis_config_tvalid = '1' else reg_poff;
      i_poff_config_reg        : process(aclk)
      begin
        if rising_edge(aclk) then
          if sclr_i = '1' then
            reg_poff <= ci_phase_adj;
          elsif aclken_i = '1' then
            reg_poff <= axi_poff_in;
          end if;
        end if;
      end process i_poff_config_reg;
    end generate i_single_channel_prog_poff;

    --Stream
    i_single_or_multi_channel_stream_poff : if C_PHASE_OFFSET = c_phase_adj_streaming generate
      axi_poff_in <= dds_poff_in;
    end generate i_single_or_multi_channel_stream_poff;

    --fixed, Multichannel
    i_mult_channel_fixed_poff : if multichannel and C_PHASE_OFFSET = c_phase_adj_fixed generate
      i_inc_ram               : dds_compiler_v5_0_lut_ram
        generic map(
          INIT_VAL     => ci_phase_adj_inits,
          C_CHANNELS   => C_CHANNELS,
          C_DATA_WIDTH => C_ACCUMULATOR_WIDTH,
          C_ADDR_WIDTH => 4,            --unnecessary, but harmless.
          C_DPRA_WIDTH => ci_chan_width,
          C_HAS_MUTE   => 1,            -- contains initial values, so mute always required
          C_HAS_CE     => 1,
          C_LATENCY    => 0
          )
        port map(
          CLK          => aclk,
          --port A
          WE           => '0',
          MUTE         => '0',          --mute_chan, REVISIT G.Old. Needs thought.
          --port B
          CE           => ce_core,
          DPRA         => std_logic_vector(master_count),
          DPO          => axi_poff_in
          );


    end generate i_mult_channel_fixed_poff;
    --Prog, Multichannel
    i_mult_channel_prog_poff : if multichannel and C_PHASE_OFFSET = c_phase_adj_prog generate
      constant ci_chan_width : integer                                          := sel_lines_reqd(C_CHANNELS);
      signal   config_poff   : std_logic_vector(C_ACCUMULATOR_WIDTH-1 downto 0) := (others => '0');
    begin
      i_poff_in_upper_tdata  : if C_PHASE_INCREMENT = c_phase_inc_prog generate
        config_poff <= s_axis_config_tdata(C_ACCUMULATOR_WIDTH + ci_byte_accum_width -1 downto ci_byte_accum_width);
      end generate i_poff_in_upper_tdata;
      i_poff_in_lower_tdata  : if C_PHASE_INCREMENT /= c_phase_inc_prog generate
        config_poff <= s_axis_config_tdata(C_ACCUMULATOR_WIDTH-1 downto 0);
      end generate i_poff_in_lower_tdata;
      i_inc_ram              : dds_compiler_v5_0_lut5_ram
        generic map(
          INIT_VAL                                                                         => ci_phase_adj_inits,
          C_CHANNELS                                                                       => C_CHANNELS,
          C_DATA_WIDTH                                                                     => C_ACCUMULATOR_WIDTH,
          C_ADDR_WIDTH                                                                     => config_write_addr'length,
          C_DPRA_WIDTH                                                                     => config_read_addr'length,
          C_HAS_MUTE                                                                       => 1,  -- contains initial values, so mute always required
          C_HAS_CE                                                                         => 1,
          C_LATENCY                                                                        => 0
          )
        port map(
          CLK                                                                              => aclk,
          --Write side
          WE                                                                               => s_axis_config_tvalid,  --REVISIT (is it necessary to
--include aclken and ready? just let the location get overwritten - the last
--write will be the valid one.
          MUTE                                                                             => '0',  --mute_chan,REVISIT - needs thought (as per if gen above)
          A                                                                                => config_write_addr,
          DI                                                                               => config_poff,
          --Read side
          CE                                                                               => ce_core,
          DPRA                                                                             => config_read_addr,  --REVISIT - needs channel addr.
          DPO                                                                              => axi_poff_in
          );

    end generate i_mult_channel_prog_poff;

  end generate i_pinc_poff_in;

  debug_interface             : if C_DEBUG_INTERFACE = 1 generate
    signal   debug_phase_nd_i : std_logic  := '0';
    constant ci_pipe          : t_pipe_top := dds_latencies.pipe;
  begin
    -- For phase validation
    debug_axi_pinc_in <= axi_pinc_in;
    debug_axi_poff_in <= axi_poff_in;
    debug_axi_chan_in <= axi_chan_in;
    debug_core_nd     <= ce_core;
    -- For sin/cos validation
    debug_phase       <= dds_debug_phase;
    i_debug_phase_in_nd_pipe  : xbip_pipe_v2_0_xst
      generic map(
        C_LATENCY  => ci_core_latency-(ci_pipe(ci_LUT_stage) +
                                      ci_pipe(ci_EFF_stage)+
                                      ci_pipe(ci_pre_op_stage)+
                                      ci_pipe(ci_op_reg_stage)),
        C_HAS_CE   => 1,
        C_HAS_SCLR => 1,
        C_WIDTH    => 1
        )
      port map(
        CLK        => aclk,
        CE         => ce_core,
        SCLR       => sclr_i,
        D(0)       => nd_i,
        Q(0)       => debug_phase_nd_i
        );
    debug_phase_nd    <= debug_phase_nd_i and ce_core;
  end generate debug_interface;

  i_dds : dds_compiler_v5_0_behv
    generic map (
      C_XDEVICEFAMILY         => C_XDEVICEFAMILY,
      C_ACCUMULATOR_WIDTH     => C_ACCUMULATOR_WIDTH,
      C_CHANNELS              => C_CHANNELS,
      C_HAS_CE                => 1,     -- always need CE to stall pipeline when FIFOs fill
      C_HAS_CHANNEL_INDEX     => boolean'pos(ci_int_core_mode.int_core = ci_int_core_mode_source),
      C_HAS_RDY               => 1,
      C_HAS_RFD               => 0,
      C_HAS_SCLR              => C_HAS_ARESETN,
      C_HAS_PHASE_OUT         => C_HAS_PHASE_OUT,
      C_HAS_PHASEGEN          => C_HAS_PHASEGEN,
      C_HAS_SINCOS            => C_HAS_SINCOS,
      C_LATENCY               => dds_pipeline_latency,  --ci_core_latency except when -1 (which is never set by GUI)
      C_MEM_TYPE              => C_MEM_TYPE,
      C_NEGATIVE_COSINE       => C_NEGATIVE_COSINE,
      C_NEGATIVE_SINE         => C_NEGATIVE_SINE,
      C_NOISE_SHAPING         => C_NOISE_SHAPING,
      C_OUTPUTS_REQUIRED      => C_OUTPUTS_REQUIRED,
      C_OUTPUT_WIDTH          => C_OUTPUT_WIDTH,
      C_PHASE_ANGLE_WIDTH     => C_PHASE_ANGLE_WIDTH,
      C_PHASE_INCREMENT       => ci_int_core_mode.phase_inc,
      C_PHASE_INCREMENT_VALUE => C_PHASE_INCREMENT_VALUE,
      C_PHASE_OFFSET          => ci_int_core_mode.phase_offset,
      C_PHASE_OFFSET_VALUE    => C_PHASE_OFFSET_VALUE,
      C_OPTIMISE_GOAL         => C_OPTIMISE_GOAL,
      C_USE_DSP48             => C_USE_DSP48,
      C_POR_MODE              => C_POR_MODE,
      C_AMPLITUDE             => C_AMPLITUDE
      )
    port map (
      ADDR                    => dds_addr,
      REG_SELECT              => dds_reg_select_dummy,
      CE                      => ce_core,
      CLK                     => aclk,
      SCLR                    => sclr_i,
      WE                      => '0',
      DATA                    => dds_data_dummy,
      PINC_IN                 => axi_pinc_in,
      POFF_IN                 => axi_poff_in,
      PHASE_IN                => axi_phase_in,
      RDY                     => dds_rdy,
      RFD                     => open,  -- always high
      CHANNEL                 => legacy_core_channel,
      COSINE                  => dds_cosine,
      SINE                    => dds_sine,
      PHASE_OUT               => dds_phase_out,
      DEBUG_PHASE             => dds_debug_phase
      );


  -----------------------------------------------------------------------------
  -- TLAST output logic
  -----------------------------------------------------------------------------

  --In this case TLAST out means 'end of TDM cycle' so is generated by the core.
  tlast_out_vector_generation : if C_HAS_TLAST = ci_tlast_vector_framing generate
    -- Pulse on last channel's output
    tlast_vector_framing      : process (aclk) is
    begin
      if rising_edge(aclk) then
        if ce_core = '1' then
          if dds_channel = std_logic_vector(to_unsigned(C_CHANNELS-2, dds_channel'length)) then
            -- get channel max one cycle earlier so that it enters the FIFO on the final channel's write
            tlast_out <= '1';
          else
            tlast_out <= '0';
          end if;
        end if;
      end if;
    end process tlast_vector_framing;
  end generate tlast_out_vector_generation;

  --FOR CONFIG TRIGGERED, see logic in CONFIG channel, as some of the required
  --signals only exist in that context.

  --In this case TLAST is completely arbitrary - just pass it through.
  tlast_out_packet_generation : if C_HAS_TLAST = ci_tlast_packet_framing generate
    axi_tlast_in <= s_phase_tlast;
  end generate tlast_out_packet_generation;

  tlast_out_diplomatic_bag : if C_HAS_TLAST = ci_tlast_packet_framing or C_HAS_TLAST = ci_tlast_config_triggered generate
    -- Propagate to output
    -- No reset required as outputs are qualified with TVALID or FIFO write enable
    tlast_delay            : xbip_pipe_v2_0_xst
      generic map(
        C_LATENCY  => dds_pipeline_latency,
        C_HAS_CE   => 1,
        C_HAS_SCLR => 0,
        C_WIDTH    => 1
        )
      port map(
        CLK        => aclk,
        CE         => ce_core,
        SCLR       => '0',
        D(0)       => axi_tlast_in,
        Q(0)       => tlast_out
        );
  end generate tlast_out_diplomatic_bag;

  -----------------------------------------------------------------------------
  -- Output channel data construction
  -----------------------------------------------------------------------------
  build_m_data_fifo_din (
    dds_cfg         => dds_cfg,
    sine            => dds_sine,
    cosine          => dds_cosine,
    channel         => dds_channel,
    user_out        => user_out,
    tlast_out       => tlast_out,
    m_data_fifo_din => m_data_fifo_din);

  build_m_phase_fifo_din (
    dds_cfg          => dds_cfg,
    phase_out        => dds_phase_out,
    channel          => dds_channel,
    user_out         => user_out,
    tlast_out        => tlast_out,
    m_phase_fifo_din => m_phase_fifo_din);

  -----------------------------------------------------------------------------
  -- Output FIFO control
  -----------------------------------------------------------------------------
  all_streaming     : if ci_int_core_mode.int_core = ci_int_core_mode_streaming generate
    no_tready       : if C_HAS_TREADY = 0 generate
      m_data_fifo_wr_enable  <= rdy_stream_i and s_axis_phase_tvalid when C_HAS_S_PHASE = 1 else rdy_stream_i;
      m_phase_fifo_wr_enable <= rdy_stream_i and s_axis_phase_tvalid when C_HAS_S_PHASE = 1 else rdy_stream_i;
    end generate no_tready;
    has_tready      : if C_HAS_TREADY = 1 generate
      m_data_fifo_wr_enable  <= rdy_stream_i and ce_core;
      m_phase_fifo_wr_enable <= rdy_stream_i and ce_core;
    end generate has_tready;
    dds_channel              <= stream_channel;
  end generate all_streaming;
  not_all_streaming : if ci_int_core_mode.int_core = ci_int_core_mode_source generate
    -- This should work for all other configurations of input channels, even if they are not present
    no_tready       : if C_HAS_TREADY = 0 generate
      m_data_fifo_wr_enable  <= dds_rdy;
      m_phase_fifo_wr_enable <= dds_rdy;
    end generate no_tready;
    has_tready      : if C_HAS_TREADY = 1 generate
      m_data_fifo_wr_enable  <= dds_rdy and ce_core;
      m_phase_fifo_wr_enable <= dds_rdy and ce_core;
    end generate has_tready;
    dds_channel              <= legacy_core_channel;
  end generate not_all_streaming;

  -----------------------------------------------------------------------------
  -- Output FIFOs
  -----------------------------------------------------------------------------

  pull_data <= m_data_fifo_not_afull and m_phase_fifo_not_afull;

  -----------------------------------------------------------------------------
  -- Set FIFO almost full threshold to one to throttle dataflow almost
  -- immediately, giving the minimum FIFO depth
  -----------------------------------------------------------------------------
  has_m_data        : if C_HAS_M_DATA = 1 generate
    i_has_tready    : if C_HAS_TREADY = 1 generate
      m_data_fifo   : glb_ifx_master_v1_0
        generic map(
          width         => m_data_fifo_width,
          depth         => m_data_fifo_depth,
          afull_thresh1 => 1,
          afull_thresh0 => 1
          )
        port map(
          aclk          => aclk,
          aclken        => aclken_i,
          areset        => sclr_i,      -- REVISIT: need to reset instantly?
          wr_enable     => m_data_fifo_wr_enable,
          wr_data       => m_data_fifo_din,
          ifx_valid     => m_axis_data_tvalid,
          ifx_ready     => m_axis_data_tready,
          ifx_data      => m_data_fifo_dout,
          full          => m_data_fifo_full,
          afull         => m_data_fifo_afull,
          not_full      => m_data_fifo_not_full,
          not_afull     => m_data_fifo_not_afull,
          add           => open
          );
    end generate i_has_tready;
    i_has_no_tready : if C_HAS_TREADY = 0 generate
      m_data_fifo_dout      <= m_data_fifo_din;
      m_axis_data_tvalid    <= m_data_fifo_wr_enable;
      m_data_fifo_not_afull <= '1';
    end generate i_has_no_tready;
  end generate has_m_data;

  has_m_phase       : if C_HAS_M_PHASE = 1 generate
    i_has_tready    : if C_HAS_TREADY = 1 generate
      m_phase_fifo  : glb_ifx_master_v1_0
        generic map(
          width         => m_phase_fifo_width,
          depth         => m_phase_fifo_depth,
          afull_thresh1 => 1,
          afull_thresh0 => 1
          )
        port map(
          aclk          => aclk,
          aclken        => aclken_i,
          areset        => sclr_i,      -- REVISIT: need to reset instantly?
          wr_enable     => m_phase_fifo_wr_enable,
          wr_data       => m_phase_fifo_din,
          ifx_valid     => m_axis_phase_tvalid,
          ifx_ready     => m_axis_phase_tready,
          ifx_data      => m_phase_fifo_dout,
          full          => m_phase_fifo_full,
          afull         => m_phase_fifo_afull,
          not_full      => m_phase_fifo_not_full,
          not_afull     => m_phase_fifo_not_afull,
          add           => open
          );
    end generate i_has_tready;
    i_has_no_tready : if C_HAS_TREADY = 0 generate
      m_phase_fifo_dout      <= m_phase_fifo_din;
      m_axis_phase_tvalid    <= m_phase_fifo_wr_enable;
      m_phase_fifo_not_afull <= '1';
    end generate i_has_no_tready;
  end generate has_m_phase;

  -----------------------------------------------------------------------------
  -- Construct output channels
  -----------------------------------------------------------------------------
  decompose_m_data_fifo_dout (
    dds_cfg           => dds_cfg,
    m_data_fifo_dout  => m_data_fifo_dout,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tlast => m_axis_data_tlast);

  decompose_m_phase_fifo_dout (
    dds_cfg            => dds_cfg,
    m_phase_fifo_dout  => m_phase_fifo_dout,
    m_axis_phase_tdata => m_axis_phase_tdata,
    m_axis_phase_tuser => m_axis_phase_tuser,
    m_axis_phase_tlast => m_axis_phase_tlast);

end architecture behavioral;
