--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:06:26 08/07/2014
-- Design Name:   
-- Module Name:   M:/vhdl/0009_00257/shift_reg/p_random_32_tb.vhd
-- Project Name:  shift_reg
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: p_random_32
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

entity p_random_32_tb is
end p_random_32_tb;

architecture behavior of p_random_32_tb is

  -- Component Declaration for the Unit Under Test (UUT)
  
  component p_random_32
    port(
      clk         : in  std_logic;
      n_reset     : in  std_logic;
      random_vect : out std_logic_vector(31 downto 0);
      ena         : in  std_logic
      );
  end component;


  --Inputs
  signal clk     : std_logic := '0';
  signal n_reset : std_logic := '0';
  signal ena     : std_logic := '0';

  --Outputs
  signal random_vect : std_logic_vector(31 downto 0);

  -- Clock period definitions
  constant clk_period : time := 10 ns;
  
begin

  -- Instantiate the Unit Under Test (UUT)
  uut : p_random_32 port map (
    clk         => clk,
    n_reset     => n_reset,
    random_vect => random_vect,
    ena         => ena
    );

  -- Clock process definitions
  clk_process : process
  begin
    clk <= '0';
    wait for clk_period/2;
    clk <= '1';
    wait for clk_period/2;
  end process;


  -- reset
  reset_proc : process
  begin
    n_reset <= '0';
    wait for 100 ns;
    n_reset <= '1';
    wait for 100 ms;
    wait;
  end process;


  -- enable process
  ena_proc : process
  begin
    ena <= '0';
    wait for 200 ns;
    wait until clk = '1';
    ena <= '1';
    wait for clk_period;
   
  end process;

  

end;
